* NGSPICE file created from multa.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

.subckt multa a[0] a[10] a[11] a[12] a[13] a[14] a[1] a[2] a[3] a[4] a[5] a[6] a[7]
+ a[8] a[9] b[0] b[10] b[11] b[12] b[13] b[14] b[15] b[16] b[17] b[18] b[1] b[2] b[3]
+ b[4] b[5] b[6] b[7] b[8] b[9] r[0] r[10] r[11] r[12] r[13] r[14] r[15] r[16] r[17]
+ r[18] r[19] r[1] r[20] r[21] r[22] r[23] r[24] r[25] r[26] r[27] r[28] r[29] r[2]
+ r[30] r[31] r[32] r[33] r[3] r[4] r[5] r[6] r[7] r[8] r[9] vccd1 vssd1
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3155_ _3731_/C vssd1 vssd1 vccd1 vccd1 _3310_/A sky130_fd_sc_hd__buf_2
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3988_ _3993_/A _3833_/B _3839_/B vssd1 vssd1 vccd1 vccd1 _3988_/Y sky130_fd_sc_hd__o21ai_1
X_5727_ _5608_/A _5608_/B _5608_/C vssd1 vssd1 vccd1 vccd1 _5727_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_10_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5658_ _5658_/A vssd1 vssd1 vccd1 vccd1 _6003_/B sky130_fd_sc_hd__buf_2
X_5589_ _5208_/B _5399_/Y _5405_/Y vssd1 vssd1 vccd1 vccd1 _5608_/A sky130_fd_sc_hd__o21ai_4
X_4609_ _4436_/Y _4442_/X _4444_/Y _4445_/X vssd1 vssd1 vccd1 vccd1 _4609_/X sky130_fd_sc_hd__o211a_1
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4960_ _4955_/Y _4957_/X _4959_/Y vssd1 vssd1 vccd1 vccd1 _4960_/Y sky130_fd_sc_hd__o21ai_1
X_3911_ _3911_/A _3911_/B _3911_/C vssd1 vssd1 vccd1 vccd1 _3912_/A sky130_fd_sc_hd__nand3_1
X_4891_ _4891_/A _4891_/B vssd1 vssd1 vccd1 vccd1 _4891_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3842_ _3821_/X _3823_/Y _3833_/X vssd1 vssd1 vccd1 vccd1 _3844_/B sky130_fd_sc_hd__o21bai_1
XFILLER_32_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5512_ _5514_/A _5514_/B _5514_/C _5643_/A vssd1 vssd1 vccd1 vccd1 _5515_/A sky130_fd_sc_hd__a22o_1
X_3773_ _5245_/A _4693_/A vssd1 vssd1 vccd1 vccd1 _3773_/Y sky130_fd_sc_hd__nand2_1
X_5443_ _5805_/A _5794_/B vssd1 vssd1 vccd1 vccd1 _5445_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5374_ _5374_/A _5378_/B vssd1 vssd1 vccd1 vccd1 _5375_/B sky130_fd_sc_hd__nand2_1
X_4325_ _4043_/C _4043_/A _4043_/B _4054_/X vssd1 vssd1 vccd1 vccd1 _4331_/B sky130_fd_sc_hd__a31oi_4
XFILLER_86_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4256_ _4251_/Y _4254_/Y _4460_/A _4255_/Y vssd1 vssd1 vccd1 vccd1 _4298_/A sky130_fd_sc_hd__o2bb2ai_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3207_ input7/X vssd1 vssd1 vccd1 vccd1 _4738_/A sky130_fd_sc_hd__clkbuf_4
X_4187_ _5123_/B vssd1 vssd1 vccd1 vccd1 _4530_/C sky130_fd_sc_hd__buf_2
X_3138_ _3521_/A vssd1 vssd1 vccd1 vccd1 _4042_/B sky130_fd_sc_hd__clkbuf_4
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4110_ _4958_/A _4110_/B vssd1 vssd1 vccd1 vccd1 _4110_/Y sky130_fd_sc_hd__nand2_2
X_5090_ _5095_/A _5095_/B _5078_/Y _5080_/X vssd1 vssd1 vccd1 vccd1 _5096_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4041_ _4041_/A vssd1 vssd1 vccd1 vccd1 _4048_/C sky130_fd_sc_hd__buf_2
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5992_ _5992_/A _5992_/B vssd1 vssd1 vccd1 vccd1 _5992_/Y sky130_fd_sc_hd__nand2_1
X_4943_ _4943_/A _4943_/B _4943_/C vssd1 vssd1 vccd1 vccd1 _4943_/X sky130_fd_sc_hd__and3_2
X_4874_ _4874_/A _4877_/D vssd1 vssd1 vccd1 vccd1 _4875_/B sky130_fd_sc_hd__nand2_2
X_3825_ input2/X vssd1 vssd1 vccd1 vccd1 _5119_/D sky130_fd_sc_hd__buf_2
X_3756_ _3761_/A _3761_/B _3756_/C vssd1 vssd1 vccd1 vccd1 _3810_/B sky130_fd_sc_hd__nand3_1
X_5426_ _5419_/Y _5420_/X _5490_/D _5490_/B vssd1 vssd1 vccd1 vccd1 _5426_/Y sky130_fd_sc_hd__o211ai_1
X_3687_ _3687_/A _3720_/C vssd1 vssd1 vccd1 vccd1 _3705_/A sky130_fd_sc_hd__or2_1
X_5357_ _5185_/X _5356_/Y _5182_/A vssd1 vssd1 vccd1 vccd1 _5519_/A sky130_fd_sc_hd__o21ai_1
XFILLER_87_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5288_ _5532_/A _5288_/B vssd1 vssd1 vccd1 vccd1 _5288_/Y sky130_fd_sc_hd__nand2_1
X_4308_ _4308_/A _4308_/B _4308_/C _4308_/D vssd1 vssd1 vccd1 vccd1 _4309_/C sky130_fd_sc_hd__nand4_1
X_4239_ _4239_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4240_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3610_ _3736_/A _3736_/B _3736_/C _3582_/C vssd1 vssd1 vccd1 vccd1 _3610_/Y sky130_fd_sc_hd__a31oi_2
X_4590_ _4877_/B _4590_/B vssd1 vssd1 vccd1 vccd1 _4751_/A sky130_fd_sc_hd__nand2_1
X_3541_ _4744_/A vssd1 vssd1 vccd1 vccd1 _4277_/C sky130_fd_sc_hd__buf_4
X_6260_ _6260_/A _6260_/B _6258_/C vssd1 vssd1 vccd1 vccd1 _6260_/X sky130_fd_sc_hd__or3b_1
X_3472_ _3472_/A _3472_/B vssd1 vssd1 vccd1 vccd1 _3478_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6191_ _6224_/A _6190_/X vssd1 vssd1 vccd1 vccd1 _6197_/A sky130_fd_sc_hd__or2b_2
X_5211_ _5211_/A _5211_/B vssd1 vssd1 vccd1 vccd1 _5403_/A sky130_fd_sc_hd__nand2_2
X_5142_ _5140_/Y _5141_/X _5126_/Y _5131_/A vssd1 vssd1 vccd1 vccd1 _5142_/X sky130_fd_sc_hd__o211a_1
X_5073_ _4751_/B _5067_/A _4885_/B _4885_/A vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__o211ai_1
XFILLER_56_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4024_ _4542_/A _4038_/B _4020_/Y _4023_/Y vssd1 vssd1 vccd1 vccd1 _4177_/A sky130_fd_sc_hd__a22o_1
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5975_ _5975_/A _5975_/B vssd1 vssd1 vccd1 vccd1 _5980_/C sky130_fd_sc_hd__nor2_2
X_4926_ _4765_/B _4924_/Y _4925_/Y vssd1 vssd1 vccd1 vccd1 _4972_/C sky130_fd_sc_hd__o21ai_2
X_4857_ _5087_/A _5087_/B _3189_/A _5376_/A vssd1 vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__o2bb2ai_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3808_ _3808_/A _3808_/B vssd1 vssd1 vccd1 vccd1 _3822_/A sky130_fd_sc_hd__nor2_1
X_4788_ _4788_/A _5530_/A _5575_/A vssd1 vssd1 vccd1 vccd1 _4788_/X sky130_fd_sc_hd__and3_1
X_3739_ _3606_/Y _3607_/Y _3856_/B _3856_/A vssd1 vssd1 vccd1 vccd1 _3739_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_79_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5409_ _3634_/X _5407_/Y _5408_/Y _5402_/Y vssd1 vssd1 vccd1 vccd1 _5413_/B sky130_fd_sc_hd__o211ai_4
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5760_ _5749_/Y _5748_/X _5751_/Y _5759_/Y _5745_/X vssd1 vssd1 vccd1 vccd1 _5761_/C
+ sky130_fd_sc_hd__o2111ai_4
X_5691_ _5673_/A _5673_/B _5690_/X vssd1 vssd1 vccd1 vccd1 _5691_/Y sky130_fd_sc_hd__a21oi_1
X_4711_ _4711_/A _4711_/B _4711_/C _4711_/D vssd1 vssd1 vccd1 vccd1 _4711_/Y sky130_fd_sc_hd__nor4_2
X_4642_ _4466_/C _4640_/Y _4641_/Y vssd1 vssd1 vccd1 vccd1 _4645_/A sky130_fd_sc_hd__o21ai_1
X_4573_ _4573_/A vssd1 vssd1 vccd1 vccd1 _4576_/A sky130_fd_sc_hd__buf_2
X_3524_ _4935_/B vssd1 vssd1 vccd1 vccd1 _4236_/B sky130_fd_sc_hd__buf_2
XFILLER_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6243_ _6244_/A _6244_/B _6244_/C vssd1 vssd1 vccd1 vccd1 _6266_/A sky130_fd_sc_hd__a21o_1
X_3455_ _4228_/A vssd1 vssd1 vccd1 vccd1 _5132_/B sky130_fd_sc_hd__buf_4
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6174_ _6173_/A _6199_/A _6173_/C _6173_/D vssd1 vssd1 vccd1 vccd1 _6240_/B sky130_fd_sc_hd__a22o_1
X_3386_ _3199_/C _3236_/Y _3312_/A vssd1 vssd1 vccd1 vccd1 _3392_/D sky130_fd_sc_hd__o21ai_2
XFILLER_69_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5125_ _5128_/A _5128_/B _5120_/A vssd1 vssd1 vccd1 vccd1 _5125_/X sky130_fd_sc_hd__a21o_1
XFILLER_29_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5056_ _5082_/A _5082_/B _5056_/C vssd1 vssd1 vccd1 vccd1 _5095_/A sky130_fd_sc_hd__nand3_2
XFILLER_84_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4007_ _3976_/A _3976_/B _3976_/C _4160_/C vssd1 vssd1 vccd1 vccd1 _4007_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_25_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5958_ _5957_/A _5957_/B _5957_/C _5957_/D vssd1 vssd1 vccd1 vccd1 _5959_/C sky130_fd_sc_hd__a22o_1
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4909_ _4913_/B _4913_/C vssd1 vssd1 vccd1 vccd1 _4909_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5889_ _5892_/A _5892_/B _5892_/C vssd1 vssd1 vccd1 vccd1 _5891_/B sky130_fd_sc_hd__nand3_1
XFILLER_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_5 _5678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3240_/A _3240_/B _3240_/C vssd1 vssd1 vccd1 vccd1 _3241_/B sky130_fd_sc_hd__nand3_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _6297_/A _3171_/B vssd1 vssd1 vccd1 vccd1 _3171_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5812_ _5808_/Y _5809_/Y _5712_/A _4829_/A _5811_/Y vssd1 vssd1 vccd1 vccd1 _5812_/X
+ sky130_fd_sc_hd__o2111a_1
X_5743_ _5743_/A vssd1 vssd1 vccd1 vccd1 _5786_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5674_ _5674_/A _5674_/B vssd1 vssd1 vccd1 vccd1 _5674_/X sky130_fd_sc_hd__or2_1
X_4625_ _4625_/A _5582_/A vssd1 vssd1 vccd1 vccd1 _4625_/Y sky130_fd_sc_hd__nand2_1
X_4556_ _4545_/A _4557_/A _4689_/A vssd1 vssd1 vccd1 vccd1 _4559_/B sky130_fd_sc_hd__nand3b_2
X_3507_ _3795_/B vssd1 vssd1 vccd1 vccd1 _4422_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4487_ _4302_/D _4486_/Y _4249_/Y vssd1 vssd1 vccd1 vccd1 _4487_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6226_ _6190_/X _6215_/Y _6224_/B vssd1 vssd1 vccd1 vccd1 _6226_/X sky130_fd_sc_hd__a21o_1
X_3438_ _3867_/A vssd1 vssd1 vccd1 vccd1 _5132_/A sky130_fd_sc_hd__clkbuf_4
X_6157_ _6156_/B _6156_/C _6156_/A vssd1 vssd1 vccd1 vccd1 _6157_/X sky130_fd_sc_hd__a21o_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _4355_/A _4366_/A _3677_/A _4235_/B vssd1 vssd1 vccd1 vccd1 _3369_/Y sky130_fd_sc_hd__nand4_4
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5310_/A _5309_/A _5309_/B vssd1 vssd1 vccd1 vccd1 _5110_/A sky130_fd_sc_hd__a21o_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ _6089_/C _6089_/B _6089_/A vssd1 vssd1 vccd1 vccd1 _6090_/A sky130_fd_sc_hd__a21o_1
X_5039_ _5035_/Y _5041_/B _5042_/A vssd1 vssd1 vccd1 vccd1 _5039_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput42 _4849_/X vssd1 vssd1 vccd1 vccd1 r[16] sky130_fd_sc_hd__buf_2
Xoutput64 _3317_/Y vssd1 vssd1 vccd1 vccd1 r[5] sky130_fd_sc_hd__buf_2
Xoutput53 _6118_/X vssd1 vssd1 vccd1 vccd1 r[26] sky130_fd_sc_hd__buf_2
XFILLER_48_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4410_ _5655_/A _4619_/B _4423_/A _4904_/B vssd1 vssd1 vccd1 vccd1 _4410_/Y sky130_fd_sc_hd__nand4_1
X_5390_ _5390_/A _6202_/B vssd1 vssd1 vccd1 vccd1 _5391_/B sky130_fd_sc_hd__nor2_1
X_4341_ _4338_/Y _4339_/X _4340_/Y _4520_/B vssd1 vssd1 vccd1 vccd1 _4341_/X sky130_fd_sc_hd__o211a_1
X_4272_ _4272_/A vssd1 vssd1 vccd1 vccd1 _4298_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3223_ _4355_/A _3223_/B vssd1 vssd1 vccd1 vccd1 _3223_/Y sky130_fd_sc_hd__nand2_1
X_6011_ _6127_/A _6127_/B _6071_/A _6065_/C _6010_/Y vssd1 vssd1 vccd1 vccd1 _6011_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_39_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3154_ _3966_/A vssd1 vssd1 vccd1 vccd1 _3731_/C sky130_fd_sc_hd__buf_2
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3987_ _3782_/X _3817_/Y _3837_/A vssd1 vssd1 vccd1 vccd1 _3987_/X sky130_fd_sc_hd__o21a_1
XFILLER_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5726_ _5726_/A vssd1 vssd1 vccd1 vccd1 _5726_/Y sky130_fd_sc_hd__inv_2
X_5657_ _5674_/B _5662_/B _5656_/Y vssd1 vssd1 vccd1 vccd1 _5657_/Y sky130_fd_sc_hd__o21ai_1
X_5588_ _5588_/A _5588_/B _5588_/C vssd1 vssd1 vccd1 vccd1 _5608_/C sky130_fd_sc_hd__nand3_4
X_4608_ _4795_/B vssd1 vssd1 vccd1 vccd1 _4643_/A sky130_fd_sc_hd__buf_2
X_4539_ _4539_/A vssd1 vssd1 vccd1 vccd1 _4832_/A sky130_fd_sc_hd__clkbuf_2
X_6209_ _6257_/B _6257_/C vssd1 vssd1 vccd1 vccd1 _6227_/A sky130_fd_sc_hd__xnor2_1
XFILLER_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3910_ _3758_/Y _3760_/Y _3755_/B vssd1 vssd1 vccd1 vccd1 _3911_/C sky130_fd_sc_hd__o21ai_2
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4890_ _4890_/A _4890_/B _4890_/C _5810_/A vssd1 vssd1 vccd1 vccd1 _4891_/B sky130_fd_sc_hd__nand4_1
X_3841_ _3835_/A _3835_/B _3836_/A vssd1 vssd1 vccd1 vccd1 _3844_/A sky130_fd_sc_hd__a21boi_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3772_ _3772_/A vssd1 vssd1 vccd1 vccd1 _5245_/A sky130_fd_sc_hd__clkbuf_4
X_5511_ _5511_/A _6283_/C _5511_/C _5514_/A vssd1 vssd1 vccd1 vccd1 _5514_/B sky130_fd_sc_hd__nand4_2
XFILLER_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5442_ _5917_/A _5808_/A _5442_/C _5810_/A vssd1 vssd1 vccd1 vccd1 _5442_/Y sky130_fd_sc_hd__nand4_2
X_5373_ _5373_/A _5658_/A vssd1 vssd1 vccd1 vccd1 _5375_/A sky130_fd_sc_hd__nand2_1
X_4324_ _4330_/B vssd1 vssd1 vccd1 vccd1 _4333_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4255_ _5119_/A vssd1 vssd1 vccd1 vccd1 _4255_/Y sky130_fd_sc_hd__inv_2
X_3206_ _3204_/Y _3205_/Y _3184_/D vssd1 vssd1 vccd1 vccd1 _3230_/C sky130_fd_sc_hd__o21ai_1
X_4186_ _4186_/A _4186_/B vssd1 vssd1 vccd1 vccd1 _4186_/Y sky130_fd_sc_hd__nand2_1
X_3137_ _4390_/A vssd1 vssd1 vccd1 vccd1 _3521_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5709_ _5799_/B _5706_/Y _5707_/Y _5708_/X vssd1 vssd1 vccd1 vccd1 _5726_/A sky130_fd_sc_hd__o211ai_2
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4040_ _3966_/A _6203_/A _4048_/B _4041_/A vssd1 vssd1 vccd1 vccd1 _4043_/A sky130_fd_sc_hd__a22o_2
XFILLER_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5991_ _5911_/A _5911_/B _5868_/C _5868_/A _5868_/B vssd1 vssd1 vccd1 vccd1 _5992_/B
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4942_ _4943_/B _4943_/C _4943_/A vssd1 vssd1 vccd1 vccd1 _4942_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4873_ _4873_/A _4873_/B vssd1 vssd1 vccd1 vccd1 _4875_/A sky130_fd_sc_hd__nand2_2
X_3824_ _3639_/X _3641_/X _3625_/Y vssd1 vssd1 vccd1 vccd1 _3824_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_32_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3755_ _3755_/A _3755_/B _3755_/C vssd1 vssd1 vccd1 vccd1 _3756_/C sky130_fd_sc_hd__nand3_1
XFILLER_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3686_ _3689_/A _3699_/A _3699_/B vssd1 vssd1 vccd1 vccd1 _3720_/C sky130_fd_sc_hd__nand3_2
X_5425_ _5427_/A _5427_/B _5256_/A _5424_/Y vssd1 vssd1 vccd1 vccd1 _5490_/B sky130_fd_sc_hd__o2bb2ai_1
X_5356_ _5172_/B _5172_/C _5172_/A vssd1 vssd1 vccd1 vccd1 _5356_/Y sky130_fd_sc_hd__a21oi_2
X_5287_ _5287_/A _5291_/A vssd1 vssd1 vccd1 vccd1 _5296_/A sky130_fd_sc_hd__nand2_1
X_4307_ _4308_/A _4308_/B _4249_/Y _4250_/X vssd1 vssd1 vccd1 vccd1 _4309_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_87_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4238_ _5299_/A _4788_/A _4238_/C _4238_/D vssd1 vssd1 vccd1 vccd1 _4238_/Y sky130_fd_sc_hd__nand4_4
X_4169_ _4166_/A _4166_/B _4520_/A _4164_/Y vssd1 vssd1 vccd1 vccd1 _4169_/X sky130_fd_sc_hd__a31o_1
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3540_ _3540_/A vssd1 vssd1 vccd1 vccd1 _3558_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3471_ _3471_/A _3471_/B vssd1 vssd1 vccd1 vccd1 _3472_/B sky130_fd_sc_hd__nor2_1
X_5210_ _3795_/B _5704_/A _5208_/Y _5209_/Y vssd1 vssd1 vccd1 vccd1 _5210_/Y sky130_fd_sc_hd__a22oi_1
X_6190_ _6190_/A _6214_/A _6190_/C vssd1 vssd1 vccd1 vccd1 _6190_/X sky130_fd_sc_hd__or3_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5141_ _5141_/A _5141_/B _5141_/C vssd1 vssd1 vccd1 vccd1 _5141_/X sky130_fd_sc_hd__and3_2
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5072_ _5095_/A _5095_/B _5070_/X _5071_/Y vssd1 vssd1 vccd1 vccd1 _5084_/A sky130_fd_sc_hd__o2bb2ai_1
X_4023_ _4540_/A _4708_/A _5696_/A _5701_/A vssd1 vssd1 vccd1 vccd1 _4023_/Y sky130_fd_sc_hd__nand4_2
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5974_ _5974_/A _5974_/B _5974_/C _5974_/D vssd1 vssd1 vccd1 vccd1 _5975_/B sky130_fd_sc_hd__nand4_1
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4925_ _4796_/A _4796_/B _4766_/A vssd1 vssd1 vccd1 vccd1 _4925_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_60_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4856_ _4863_/A vssd1 vssd1 vccd1 vccd1 _5376_/A sky130_fd_sc_hd__inv_2
X_3807_ _3803_/X _3806_/X _3799_/Y _3793_/Y vssd1 vssd1 vccd1 vccd1 _3808_/B sky130_fd_sc_hd__o211a_1
XFILLER_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4787_ _5037_/B vssd1 vssd1 vccd1 vccd1 _5449_/A sky130_fd_sc_hd__clkbuf_4
X_3738_ _3736_/X _3737_/Y _3733_/Y _3734_/X vssd1 vssd1 vccd1 vccd1 _3856_/A sky130_fd_sc_hd__o211a_1
X_3669_ _3669_/A vssd1 vssd1 vccd1 vccd1 _3669_/X sky130_fd_sc_hd__clkbuf_8
X_5408_ _5248_/Y _5263_/B _5244_/Y vssd1 vssd1 vccd1 vccd1 _5408_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_87_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5339_ _5339_/A _5339_/B _5339_/C vssd1 vssd1 vccd1 vccd1 _5351_/A sky130_fd_sc_hd__nand3_2
XFILLER_87_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5690_ _5654_/A _6137_/C _5852_/C _5652_/X vssd1 vssd1 vccd1 vccd1 _5690_/X sky130_fd_sc_hd__a31o_1
XFILLER_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4710_ _4711_/A _4711_/C _4711_/D _4711_/B vssd1 vssd1 vccd1 vccd1 _4710_/X sky130_fd_sc_hd__o22a_1
X_4641_ _4641_/A _4641_/B vssd1 vssd1 vccd1 vccd1 _4641_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4572_ _5231_/A _4753_/D vssd1 vssd1 vccd1 vccd1 _4573_/A sky130_fd_sc_hd__nand2_1
X_3523_ _3465_/Y _3446_/X _3452_/Y vssd1 vssd1 vccd1 vccd1 _3561_/A sky130_fd_sc_hd__a21boi_1
X_6242_ _6257_/A _6242_/B vssd1 vssd1 vccd1 vccd1 _6244_/C sky130_fd_sc_hd__xor2_1
X_3454_ _3376_/Y _3372_/B _3360_/A vssd1 vssd1 vccd1 vccd1 _3574_/B sky130_fd_sc_hd__a21boi_1
X_6173_ _6173_/A _6199_/A _6173_/C _6173_/D vssd1 vssd1 vccd1 vccd1 _6240_/C sky130_fd_sc_hd__nand4_2
X_3385_ _3483_/A _3484_/A _3384_/X vssd1 vssd1 vccd1 vccd1 _3388_/B sky130_fd_sc_hd__a21o_1
X_5124_ _5124_/A _5124_/B vssd1 vssd1 vccd1 vccd1 _5128_/A sky130_fd_sc_hd__nand2_2
X_5055_ _4853_/B _5232_/A _3223_/B _5372_/C _5081_/A vssd1 vssd1 vccd1 vccd1 _5056_/C
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_84_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4006_ _3976_/B _3976_/C _3976_/A vssd1 vssd1 vccd1 vccd1 _4006_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_25_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5957_ _5957_/A _5957_/B _5957_/C _5957_/D vssd1 vssd1 vccd1 vccd1 _5959_/B sky130_fd_sc_hd__nand4_1
X_4908_ _4776_/B _4907_/X _5656_/A _5534_/A _4903_/Y vssd1 vssd1 vccd1 vccd1 _4913_/C
+ sky130_fd_sc_hd__o2111ai_2
X_5888_ _5884_/Y _5885_/Y _5886_/X _5887_/Y vssd1 vssd1 vccd1 vccd1 _5892_/C sky130_fd_sc_hd__o22ai_4
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4839_ _4839_/A _4839_/B _4839_/C vssd1 vssd1 vccd1 vccd1 _4845_/B sky130_fd_sc_hd__nand3_2
XFILLER_88_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_6 _5678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _3170_/A _3170_/B vssd1 vssd1 vccd1 vccd1 _3171_/B sky130_fd_sc_hd__nor2_2
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5811_ _5811_/A _5811_/B vssd1 vssd1 vccd1 vccd1 _5811_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5742_ _5673_/Y _5675_/X _5741_/Y vssd1 vssd1 vccd1 vccd1 _5742_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5673_ _5673_/A _5673_/B vssd1 vssd1 vccd1 vccd1 _5673_/Y sky130_fd_sc_hd__nand2_2
X_4624_ _4257_/Y _4473_/X _4456_/B _4458_/Y vssd1 vssd1 vccd1 vccd1 _4628_/A sky130_fd_sc_hd__a22o_1
X_4555_ _4414_/X _4550_/X _4420_/X vssd1 vssd1 vccd1 vccd1 _4559_/A sky130_fd_sc_hd__a21bo_1
X_3506_ _5037_/A vssd1 vssd1 vccd1 vccd1 _3795_/B sky130_fd_sc_hd__buf_4
X_4486_ _4237_/X _4241_/X _4381_/Y _4382_/X vssd1 vssd1 vccd1 vccd1 _4486_/Y sky130_fd_sc_hd__a31oi_1
X_6225_ _6195_/Y _6221_/Y _6274_/A vssd1 vssd1 vccd1 vccd1 _6225_/Y sky130_fd_sc_hd__o21bai_1
X_3437_ _3437_/A vssd1 vssd1 vccd1 vccd1 _3867_/A sky130_fd_sc_hd__buf_2
X_6156_ _6156_/A _6156_/B _6156_/C vssd1 vssd1 vccd1 vccd1 _6156_/Y sky130_fd_sc_hd__nand3_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _3368_/A _3368_/B vssd1 vssd1 vccd1 vccd1 _3368_/Y sky130_fd_sc_hd__nand2_1
X_5107_ _5107_/A vssd1 vssd1 vccd1 vccd1 _5325_/A sky130_fd_sc_hd__clkbuf_2
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6087_ _6087_/A _6087_/B vssd1 vssd1 vccd1 vccd1 _6089_/A sky130_fd_sc_hd__nand2_1
X_3299_ _3293_/Y _3226_/A _3296_/Y _3298_/X vssd1 vssd1 vccd1 vccd1 _3300_/D sky130_fd_sc_hd__o211ai_2
XFILLER_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5038_ _4903_/A _4902_/A _4904_/Y _5037_/Y vssd1 vssd1 vccd1 vccd1 _5042_/A sky130_fd_sc_hd__a22oi_2
XFILLER_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput43 _5018_/X vssd1 vssd1 vccd1 vccd1 r[17] sky130_fd_sc_hd__buf_2
Xoutput54 _6163_/X vssd1 vssd1 vccd1 vccd1 r[27] sky130_fd_sc_hd__buf_2
Xoutput65 _3397_/X vssd1 vssd1 vccd1 vccd1 r[6] sky130_fd_sc_hd__buf_2
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4340_ _4340_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4340_/Y sky130_fd_sc_hd__nand2_1
X_4271_ _4063_/Y _4259_/X _4266_/Y _4270_/Y vssd1 vssd1 vccd1 vccd1 _4272_/A sky130_fd_sc_hd__o211ai_1
X_6010_ _6010_/A _6010_/B vssd1 vssd1 vccd1 vccd1 _6010_/Y sky130_fd_sc_hd__nand2_1
X_3222_ _5231_/A vssd1 vssd1 vccd1 vccd1 _3223_/B sky130_fd_sc_hd__buf_6
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3153_ _3514_/A vssd1 vssd1 vccd1 vccd1 _3966_/A sky130_fd_sc_hd__buf_2
XFILLER_82_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3986_ _3984_/X _3985_/Y _3973_/B _3975_/B vssd1 vssd1 vccd1 vccd1 _3990_/B sky130_fd_sc_hd__o211ai_1
XFILLER_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5725_ _5729_/A _5729_/B _5728_/A vssd1 vssd1 vccd1 vccd1 _5725_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_10_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5656_ _5656_/A _5917_/C vssd1 vssd1 vccd1 vccd1 _5656_/Y sky130_fd_sc_hd__nand2_1
X_4607_ _4607_/A _4607_/B _4607_/C vssd1 vssd1 vccd1 vccd1 _4795_/B sky130_fd_sc_hd__nand3_1
X_5587_ _5571_/Y _5573_/Y _5372_/Y vssd1 vssd1 vccd1 vccd1 _5588_/C sky130_fd_sc_hd__o21ai_4
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4538_ _4956_/A _5299_/C _4384_/A _4714_/A vssd1 vssd1 vccd1 vccd1 _4539_/A sky130_fd_sc_hd__a22o_1
X_4469_ _4466_/A _4466_/B _4466_/C vssd1 vssd1 vccd1 vccd1 _4469_/Y sky130_fd_sc_hd__a21oi_2
X_6208_ _6208_/A _6208_/B vssd1 vssd1 vccd1 vccd1 _6257_/C sky130_fd_sc_hd__and2_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6139_ _6131_/X _6139_/B _6139_/C vssd1 vssd1 vccd1 vccd1 _6143_/A sky130_fd_sc_hd__nand3b_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3840_ _3847_/A _3847_/B _3847_/C vssd1 vssd1 vccd1 vccd1 _3840_/X sky130_fd_sc_hd__and3_1
X_3771_ _3418_/A _5378_/A _4532_/A _4423_/A _3770_/Y vssd1 vssd1 vccd1 vccd1 _3771_/X
+ sky130_fd_sc_hd__a41o_1
X_5510_ _5513_/A _5513_/B _5510_/C _5643_/B vssd1 vssd1 vccd1 vccd1 _5776_/A sky130_fd_sc_hd__nand4_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5441_ _5288_/Y _5296_/D _5290_/Y vssd1 vssd1 vccd1 vccd1 _5451_/A sky130_fd_sc_hd__a21oi_1
X_5372_ _5597_/A _5372_/B _5372_/C _5831_/B vssd1 vssd1 vccd1 vccd1 _5372_/Y sky130_fd_sc_hd__nand4_2
X_4323_ _4323_/A _4323_/B _4323_/C vssd1 vssd1 vccd1 vccd1 _4330_/B sky130_fd_sc_hd__nand3_1
XFILLER_86_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4254_ _4254_/A _4254_/B vssd1 vssd1 vccd1 vccd1 _4254_/Y sky130_fd_sc_hd__nand2_2
X_4185_ _4020_/B _4365_/A _3639_/A _6010_/A _4182_/Y vssd1 vssd1 vccd1 vccd1 _4213_/B
+ sky130_fd_sc_hd__o2111ai_2
X_3205_ _3791_/C _3179_/C _5006_/A _3218_/A vssd1 vssd1 vccd1 vccd1 _3205_/Y sky130_fd_sc_hd__a22oi_1
X_3136_ _4176_/A vssd1 vssd1 vccd1 vccd1 _4390_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5708_ _5799_/A _5698_/Y _5704_/Y vssd1 vssd1 vccd1 vccd1 _5708_/X sky130_fd_sc_hd__a21o_1
X_3969_ _3799_/Y _3804_/X _3793_/Y vssd1 vssd1 vccd1 vccd1 _4010_/C sky130_fd_sc_hd__a21boi_2
X_5639_ _5639_/A _5639_/B _5639_/C vssd1 vssd1 vccd1 vccd1 _5776_/C sky130_fd_sc_hd__nand3_1
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5990_ _5868_/A _5868_/B _5868_/C _5989_/Y vssd1 vssd1 vccd1 vccd1 _5992_/A sky130_fd_sc_hd__a31o_1
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4941_ _4941_/A _5718_/A vssd1 vssd1 vccd1 vccd1 _4943_/A sky130_fd_sc_hd__nand2_1
X_4872_ _5931_/A vssd1 vssd1 vccd1 vccd1 _5407_/C sky130_fd_sc_hd__buf_4
XFILLER_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3823_ _3837_/C _3837_/A _3837_/B vssd1 vssd1 vccd1 vccd1 _3823_/Y sky130_fd_sc_hd__a21oi_2
X_3754_ _3754_/A _3754_/B vssd1 vssd1 vccd1 vccd1 _3761_/B sky130_fd_sc_hd__nand2_1
X_3685_ _3685_/A _3685_/B _3685_/C vssd1 vssd1 vccd1 vccd1 _3699_/B sky130_fd_sc_hd__nand3_2
X_5424_ _5424_/A _5424_/B vssd1 vssd1 vccd1 vccd1 _5424_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5355_ _5355_/A _5355_/B _5355_/C vssd1 vssd1 vccd1 vccd1 _5520_/B sky130_fd_sc_hd__nand3_2
X_4306_ _4124_/B _4131_/Y _4124_/C vssd1 vssd1 vccd1 vccd1 _4309_/A sky130_fd_sc_hd__o21ai_1
X_5286_ _5286_/A _5286_/B vssd1 vssd1 vccd1 vccd1 _5291_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4237_ _4087_/Y _4088_/Y _4235_/Y _4236_/Y vssd1 vssd1 vccd1 vccd1 _4237_/X sky130_fd_sc_hd__a22o_2
XFILLER_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4168_ _4338_/A _4164_/Y _4167_/X vssd1 vssd1 vccd1 vccd1 _4168_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4099_ _4100_/A _4100_/B _4100_/C vssd1 vssd1 vccd1 vccd1 _4130_/A sky130_fd_sc_hd__a21oi_2
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3470_ _3419_/Y _3421_/Y _3423_/Y vssd1 vssd1 vccd1 vccd1 _3471_/B sky130_fd_sc_hd__a21oi_1
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5140_ _5141_/B _5141_/C _5141_/A vssd1 vssd1 vccd1 vccd1 _5140_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5071_ _5080_/A _5070_/C _5070_/A vssd1 vssd1 vccd1 vccd1 _5071_/Y sky130_fd_sc_hd__a21oi_1
X_4022_ _5119_/D vssd1 vssd1 vccd1 vccd1 _5701_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5973_ _5984_/A _5984_/B vssd1 vssd1 vccd1 vccd1 _6193_/A sky130_fd_sc_hd__xnor2_4
XFILLER_25_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4924_ _4924_/A _4924_/B vssd1 vssd1 vccd1 vccd1 _4924_/Y sky130_fd_sc_hd__nand2_2
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4855_ _4855_/A _4855_/B _5059_/A _5237_/A vssd1 vssd1 vccd1 vccd1 _5087_/B sky130_fd_sc_hd__nand4_2
XFILLER_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3806_ _3806_/A _5994_/B _3966_/B vssd1 vssd1 vccd1 vccd1 _3806_/X sky130_fd_sc_hd__and3_1
X_4786_ _4786_/A _4786_/B _4786_/C vssd1 vssd1 vccd1 vccd1 _4951_/A sky130_fd_sc_hd__nand3_4
X_3737_ _3609_/A _3609_/B _3609_/C _3607_/A vssd1 vssd1 vccd1 vccd1 _3737_/Y sky130_fd_sc_hd__a31oi_4
X_3668_ _3657_/A _3564_/B _3564_/A vssd1 vssd1 vccd1 vccd1 _3708_/A sky130_fd_sc_hd__a21boi_1
X_5407_ _5407_/A _5407_/B _5407_/C vssd1 vssd1 vccd1 vccd1 _5407_/Y sky130_fd_sc_hd__nand3_1
X_3599_ _3857_/B _3597_/Y _6295_/A vssd1 vssd1 vccd1 vccd1 _3600_/C sky130_fd_sc_hd__o21ai_2
X_5338_ _5150_/Y _5336_/Y _5163_/B _5337_/X _5332_/B vssd1 vssd1 vccd1 vccd1 _5339_/C
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5269_ _5269_/A _5424_/A _5424_/B vssd1 vssd1 vccd1 vccd1 _5431_/A sky130_fd_sc_hd__nand3_2
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4640_ _4640_/A _4640_/B vssd1 vssd1 vccd1 vccd1 _4640_/Y sky130_fd_sc_hd__nand2_1
X_4571_ _4571_/A _4571_/B _5065_/B _5570_/A vssd1 vssd1 vccd1 vccd1 _4576_/C sky130_fd_sc_hd__nand4_4
X_3522_ _3522_/A _5994_/A _3730_/A _3522_/D vssd1 vssd1 vccd1 vccd1 _3730_/B sky130_fd_sc_hd__nand4_4
X_6241_ _6257_/B _6257_/C _6240_/X vssd1 vssd1 vccd1 vccd1 _6242_/B sky130_fd_sc_hd__a21oi_1
X_3453_ _3465_/A _3465_/B _3446_/X _3452_/Y vssd1 vssd1 vccd1 vccd1 _3574_/A sky130_fd_sc_hd__a22o_1
XFILLER_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6172_ _6198_/A _6171_/B _5825_/D _4830_/A vssd1 vssd1 vccd1 vccd1 _6173_/D sky130_fd_sc_hd__a2bb2o_1
X_3384_ _3389_/A _3487_/A vssd1 vssd1 vccd1 vccd1 _3384_/X sky130_fd_sc_hd__or2_1
X_5123_ _5123_/A _5123_/B vssd1 vssd1 vccd1 vccd1 _5124_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _5245_/B vssd1 vssd1 vccd1 vccd1 _5372_/C sky130_fd_sc_hd__buf_4
XFILLER_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4005_ _4005_/A _4005_/B vssd1 vssd1 vccd1 vccd1 _4005_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_25_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5956_ _5956_/A _5956_/B vssd1 vssd1 vccd1 vccd1 _5957_/D sky130_fd_sc_hd__nand2_1
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5887_ _5872_/Y _5879_/Y _5881_/X vssd1 vssd1 vccd1 vccd1 _5887_/Y sky130_fd_sc_hd__a21boi_1
X_4907_ _5025_/A vssd1 vssd1 vccd1 vccd1 _4907_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4838_ _4827_/X _4832_/X _4824_/Y _4819_/Y vssd1 vssd1 vccd1 vccd1 _4839_/C sky130_fd_sc_hd__o211ai_1
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4769_ _4576_/A _4579_/Y _4576_/C _4745_/Y vssd1 vssd1 vccd1 vccd1 _4769_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_20_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_7 _3150_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5810_ _5810_/A _5810_/B vssd1 vssd1 vccd1 vccd1 _5811_/A sky130_fd_sc_hd__nand2_2
X_5741_ _5673_/Y _5675_/X _5684_/Y vssd1 vssd1 vccd1 vccd1 _5741_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5672_ _5652_/X _5654_/X _5673_/B _5673_/A vssd1 vssd1 vccd1 vccd1 _5672_/X sky130_fd_sc_hd__o211a_4
X_4623_ _4623_/A _4623_/B _4623_/C vssd1 vssd1 vccd1 vccd1 _4635_/A sky130_fd_sc_hd__nand3_4
X_4554_ _4546_/Y _4549_/X _4551_/Y _4553_/X vssd1 vssd1 vccd1 vccd1 _4554_/Y sky130_fd_sc_hd__o211ai_4
X_3505_ _5212_/A vssd1 vssd1 vccd1 vccd1 _5037_/A sky130_fd_sc_hd__clkbuf_2
X_6224_ _6224_/A _6224_/B _6223_/X vssd1 vssd1 vccd1 vccd1 _6274_/A sky130_fd_sc_hd__or3b_2
X_4485_ _4489_/C _4467_/A _4641_/A vssd1 vssd1 vccd1 vccd1 _4490_/A sky130_fd_sc_hd__a21o_1
X_3436_ _3429_/Y _3433_/Y _3342_/B _3530_/A vssd1 vssd1 vccd1 vccd1 _3439_/A sky130_fd_sc_hd__o2bb2ai_2
X_6155_ _6104_/B _6123_/X _6153_/Y vssd1 vssd1 vccd1 vccd1 _6156_/C sky130_fd_sc_hd__a21o_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _3368_/A _3368_/B _3366_/Y vssd1 vssd1 vccd1 vccd1 _3367_/Y sky130_fd_sc_hd__o21ai_2
X_6086_ _6143_/C _6061_/X _6083_/Y _6085_/X vssd1 vssd1 vccd1 vccd1 _6094_/B sky130_fd_sc_hd__o211ai_2
X_5106_ _5278_/B _5098_/Y _5103_/Y _5105_/X vssd1 vssd1 vccd1 vccd1 _5107_/A sky130_fd_sc_hd__o211ai_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3298_ _3345_/B _3287_/X _3345_/A vssd1 vssd1 vccd1 vccd1 _3298_/X sky130_fd_sc_hd__a21o_1
X_5037_ _5037_/A _5037_/B vssd1 vssd1 vccd1 vccd1 _5037_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5939_ _5848_/Y _5855_/X _5840_/Y vssd1 vssd1 vccd1 vccd1 _5940_/C sky130_fd_sc_hd__a21boi_2
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput66 _6295_/X vssd1 vssd1 vccd1 vccd1 r[7] sky130_fd_sc_hd__buf_2
Xoutput44 _5197_/X vssd1 vssd1 vccd1 vccd1 r[18] sky130_fd_sc_hd__buf_2
Xoutput55 _6197_/X vssd1 vssd1 vccd1 vccd1 r[28] sky130_fd_sc_hd__buf_2
XFILLER_95_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4270_ _4270_/A _4761_/B _4277_/C vssd1 vssd1 vccd1 vccd1 _4270_/Y sky130_fd_sc_hd__nand3_2
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3221_ _3908_/A vssd1 vssd1 vccd1 vccd1 _5231_/A sky130_fd_sc_hd__buf_4
XFILLER_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3152_ _4176_/A vssd1 vssd1 vccd1 vccd1 _3514_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3985_ _3985_/A _3985_/B vssd1 vssd1 vccd1 vccd1 _3985_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5724_ _5724_/A vssd1 vssd1 vccd1 vccd1 _5728_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5655_ _5655_/A _5658_/A vssd1 vssd1 vccd1 vccd1 _5662_/B sky130_fd_sc_hd__nand2_2
X_4606_ _4599_/B _4606_/B _4606_/C vssd1 vssd1 vccd1 vccd1 _4607_/C sky130_fd_sc_hd__nand3b_1
X_5586_ _5674_/A _5674_/B _5583_/B _5654_/A vssd1 vssd1 vccd1 vccd1 _5588_/B sky130_fd_sc_hd__o211ai_4
X_4537_ _4557_/B vssd1 vssd1 vccd1 vccd1 _4689_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4468_ _4468_/A _4641_/B vssd1 vssd1 vccd1 vccd1 _4468_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6207_ _6205_/C _6236_/C _6253_/A _6206_/B _6244_/B vssd1 vssd1 vccd1 vccd1 _6208_/B
+ sky130_fd_sc_hd__a32o_1
X_3419_ _3419_/A _3419_/B vssd1 vssd1 vccd1 vccd1 _3419_/Y sky130_fd_sc_hd__nand2_2
X_6138_ _6138_/A _6138_/B vssd1 vssd1 vccd1 vccd1 _6139_/C sky130_fd_sc_hd__nor2_1
X_4399_ _4399_/A _4399_/B vssd1 vssd1 vccd1 vccd1 _4400_/C sky130_fd_sc_hd__nor2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6069_ _6010_/Y _6012_/Y _6006_/D vssd1 vssd1 vccd1 vccd1 _6069_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_26_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3770_ _4369_/A _4884_/A vssd1 vssd1 vccd1 vccd1 _3770_/Y sky130_fd_sc_hd__nand2_2
X_5440_ _5464_/A _5465_/A _4417_/X _6171_/C vssd1 vssd1 vccd1 vccd1 _5460_/B sky130_fd_sc_hd__a211o_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5371_ _5236_/B _5236_/A _5420_/C _5420_/B vssd1 vssd1 vccd1 vccd1 _5371_/Y sky130_fd_sc_hd__a22oi_2
X_4322_ _4322_/A _4322_/B _4322_/C vssd1 vssd1 vccd1 vccd1 _4323_/C sky130_fd_sc_hd__nand3_1
X_4253_ _4874_/A _5286_/B vssd1 vssd1 vccd1 vccd1 _4254_/B sky130_fd_sc_hd__nand2_1
X_3204_ _3639_/B _3204_/B vssd1 vssd1 vccd1 vccd1 _3204_/Y sky130_fd_sc_hd__nand2_1
X_4184_ _4184_/A _5284_/D vssd1 vssd1 vccd1 vccd1 _4365_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3135_ _3218_/A vssd1 vssd1 vccd1 vccd1 _3190_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3968_ _3968_/A _4143_/A _4143_/B vssd1 vssd1 vccd1 vccd1 _4052_/A sky130_fd_sc_hd__nor3_2
XFILLER_23_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5707_ _5538_/X _5540_/X _5554_/B _5542_/Y vssd1 vssd1 vccd1 vccd1 _5707_/Y sky130_fd_sc_hd__a2bb2oi_1
X_3899_ _4874_/A _4930_/A vssd1 vssd1 vccd1 vccd1 _3902_/B sky130_fd_sc_hd__nand2_2
X_5638_ _5638_/A _5640_/C _5640_/D vssd1 vssd1 vccd1 vccd1 _5639_/C sky130_fd_sc_hd__nand3_1
X_5569_ _5625_/A _5625_/B vssd1 vssd1 vccd1 vccd1 _5618_/A sky130_fd_sc_hd__nand2_1
XFILLER_2_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4940_ _5132_/A _5436_/B _5434_/D _3783_/A vssd1 vssd1 vccd1 vccd1 _4943_/C sky130_fd_sc_hd__a22o_2
XFILLER_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4871_ _4871_/A vssd1 vssd1 vccd1 vccd1 _4871_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3822_ _3822_/A _3822_/B _3822_/C vssd1 vssd1 vccd1 vccd1 _3837_/C sky130_fd_sc_hd__nand3_2
X_3753_ _4744_/A _3774_/B vssd1 vssd1 vccd1 vccd1 _3754_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3684_ _3684_/A _3684_/B vssd1 vssd1 vccd1 vccd1 _3685_/C sky130_fd_sc_hd__nor2_1
X_5423_ _5430_/A _5614_/A _5423_/C _5423_/D vssd1 vssd1 vccd1 vccd1 _5490_/D sky130_fd_sc_hd__nand4_2
X_5354_ _5513_/A _5364_/A _5354_/C vssd1 vssd1 vccd1 vccd1 _5355_/C sky130_fd_sc_hd__nand3_1
X_4305_ _4131_/Y _4227_/X _4297_/Y _4304_/X vssd1 vssd1 vccd1 vccd1 _4322_/B sky130_fd_sc_hd__o211ai_4
X_5285_ _5285_/A _5448_/A vssd1 vssd1 vccd1 vccd1 _5287_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4236_ _4236_/A _4236_/B vssd1 vssd1 vccd1 vccd1 _4236_/Y sky130_fd_sc_hd__nand2_1
X_4167_ _4338_/A _4520_/B _4164_/Y vssd1 vssd1 vccd1 vccd1 _4167_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4098_ _4097_/Y _3911_/C _3927_/C vssd1 vssd1 vccd1 vccd1 _4098_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_55_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5070_ _5070_/A _5080_/A _5070_/C vssd1 vssd1 vccd1 vccd1 _5070_/X sky130_fd_sc_hd__and3_1
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4021_ _5123_/B vssd1 vssd1 vccd1 vccd1 _5696_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5972_ _5883_/A _5883_/B _5883_/C _5892_/C _5892_/A vssd1 vssd1 vccd1 vccd1 _5984_/B
+ sky130_fd_sc_hd__a32oi_4
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4923_ _4919_/Y _4922_/X _4981_/B _4981_/C vssd1 vssd1 vccd1 vccd1 _4972_/B sky130_fd_sc_hd__o211ai_2
XFILLER_33_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4854_ _5230_/A vssd1 vssd1 vccd1 vccd1 _5237_/A sky130_fd_sc_hd__buf_2
XFILLER_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3805_ _3793_/Y _3799_/Y _3804_/X vssd1 vssd1 vccd1 vccd1 _3808_/A sky130_fd_sc_hd__a21oi_2
X_4785_ _4473_/X _4592_/B _4593_/Y _4589_/Y vssd1 vssd1 vccd1 vccd1 _4786_/C sky130_fd_sc_hd__o22ai_4
X_3736_ _3736_/A _3736_/B _3736_/C vssd1 vssd1 vccd1 vccd1 _3736_/X sky130_fd_sc_hd__and3_1
X_3667_ _3685_/A vssd1 vssd1 vccd1 vccd1 _3667_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5406_ _5263_/A _5249_/Y _5402_/Y _5405_/Y vssd1 vssd1 vccd1 vccd1 _5413_/A sky130_fd_sc_hd__a22o_1
X_3598_ _3598_/A _3598_/B _3598_/C vssd1 vssd1 vccd1 vccd1 _6295_/A sky130_fd_sc_hd__nor3_4
X_5337_ _5337_/A vssd1 vssd1 vccd1 vccd1 _5337_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5268_ _5268_/A _5268_/B _5420_/B _5420_/C vssd1 vssd1 vccd1 vccd1 _5424_/B sky130_fd_sc_hd__nand4_2
X_4219_ _4219_/A _4219_/B vssd1 vssd1 vccd1 vccd1 _4220_/D sky130_fd_sc_hd__nand2_1
X_5199_ _5171_/C _5170_/B _5171_/D vssd1 vssd1 vccd1 vccd1 _5339_/A sky130_fd_sc_hd__a21boi_1
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4570_ _4863_/A vssd1 vssd1 vccd1 vccd1 _5570_/A sky130_fd_sc_hd__buf_2
X_3521_ _3521_/A _3639_/B _5850_/A vssd1 vssd1 vccd1 vccd1 _3522_/D sky130_fd_sc_hd__and3_1
XFILLER_6_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6240_ _6240_/A _6240_/B _6240_/C _6240_/D vssd1 vssd1 vccd1 vccd1 _6240_/X sky130_fd_sc_hd__and4_1
X_3452_ _3452_/A _3452_/B _3452_/C vssd1 vssd1 vccd1 vccd1 _3452_/Y sky130_fd_sc_hd__nand3_2
X_6171_ _6171_/A _6171_/B _6171_/C _6198_/A vssd1 vssd1 vccd1 vccd1 _6173_/C sky130_fd_sc_hd__or4_1
X_3383_ _3389_/A _3487_/A _3483_/A _3484_/A vssd1 vssd1 vccd1 vccd1 _3388_/A sky130_fd_sc_hd__o211ai_1
X_5122_ _4932_/A _4932_/B _4935_/Y _4936_/Y vssd1 vssd1 vccd1 vccd1 _5122_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5053_ _5053_/A _5240_/D vssd1 vssd1 vccd1 vccd1 _5232_/A sky130_fd_sc_hd__nand2_2
XFILLER_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4004_ _4004_/A _4004_/B vssd1 vssd1 vccd1 vccd1 _4005_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5955_ _5960_/B _5960_/C vssd1 vssd1 vccd1 vccd1 _5956_/B sky130_fd_sc_hd__nand2_1
X_5886_ _5748_/X _5740_/X _5872_/Y _5879_/Y vssd1 vssd1 vccd1 vccd1 _5886_/X sky130_fd_sc_hd__o211a_1
XFILLER_80_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4906_ _4906_/A _4906_/B vssd1 vssd1 vccd1 vccd1 _5025_/A sky130_fd_sc_hd__nand2_2
XFILLER_40_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4837_ _4832_/A _4687_/Y _4819_/Y _4824_/Y vssd1 vssd1 vccd1 vccd1 _4839_/B sky130_fd_sc_hd__a22o_1
X_4768_ _4746_/A _4746_/B _4745_/A vssd1 vssd1 vccd1 vccd1 _4768_/Y sky130_fd_sc_hd__a21oi_2
X_4699_ input3/X vssd1 vssd1 vccd1 vccd1 _5288_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3719_ _3719_/A _3719_/B _3719_/C vssd1 vssd1 vccd1 vccd1 _3720_/D sky130_fd_sc_hd__nand3_1
XFILLER_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_8 _6297_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5740_ _5734_/Y _5738_/Y _5739_/X _5723_/Y vssd1 vssd1 vccd1 vccd1 _5740_/X sky130_fd_sc_hd__o211a_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _5826_/A _5826_/B _5671_/C vssd1 vssd1 vccd1 vccd1 _5673_/A sky130_fd_sc_hd__nand3_2
X_4622_ _4458_/Y _4453_/Y _4456_/B vssd1 vssd1 vccd1 vccd1 _4623_/C sky130_fd_sc_hd__o21ai_1
X_4553_ _4557_/A _4689_/A _4689_/B vssd1 vssd1 vccd1 vccd1 _4553_/X sky130_fd_sc_hd__a21o_1
X_4484_ _4484_/A _4484_/B vssd1 vssd1 vccd1 vccd1 _4641_/A sky130_fd_sc_hd__nand2_2
X_3504_ _3504_/A vssd1 vssd1 vccd1 vccd1 _3641_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6223_ _6190_/C _6214_/A _6190_/A _6215_/Y vssd1 vssd1 vccd1 vccd1 _6223_/X sky130_fd_sc_hd__o31a_1
X_3435_ _4861_/A _3774_/B vssd1 vssd1 vccd1 vccd1 _3530_/A sky130_fd_sc_hd__nand2_4
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6154_ _6101_/A _6101_/B _6123_/X _6153_/Y vssd1 vssd1 vccd1 vccd1 _6156_/B sky130_fd_sc_hd__o211ai_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _4201_/A _5248_/A vssd1 vssd1 vccd1 vccd1 _3366_/Y sky130_fd_sc_hd__nand2_2
X_6085_ _6089_/C _6089_/B _6084_/Y vssd1 vssd1 vccd1 vccd1 _6085_/X sky130_fd_sc_hd__a21o_1
X_5105_ _5278_/A _5203_/A _5085_/A vssd1 vssd1 vccd1 vccd1 _5105_/X sky130_fd_sc_hd__a21o_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ _5087_/C _4366_/A vssd1 vssd1 vccd1 vccd1 _3345_/A sky130_fd_sc_hd__nand2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5034_/A _5034_/B _4903_/B _5208_/A _5025_/Y vssd1 vssd1 vccd1 vccd1 _5041_/B
+ sky130_fd_sc_hd__o221ai_4
XFILLER_38_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5938_ _5935_/A _5935_/B _5942_/C _5942_/B vssd1 vssd1 vccd1 vccd1 _5940_/B sky130_fd_sc_hd__o211ai_1
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5869_ _5673_/Y _5675_/X _5741_/Y _5860_/B vssd1 vssd1 vccd1 vccd1 _5869_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput45 _5363_/Y vssd1 vssd1 vccd1 vccd1 r[19] sky130_fd_sc_hd__buf_2
Xoutput56 _6218_/Y vssd1 vssd1 vccd1 vccd1 r[29] sky130_fd_sc_hd__buf_2
Xoutput67 _3601_/Y vssd1 vssd1 vccd1 vccd1 r[8] sky130_fd_sc_hd__buf_2
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3220_ _4025_/A vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__clkbuf_4
X_3151_ _3151_/A vssd1 vssd1 vccd1 vccd1 _6297_/A sky130_fd_sc_hd__buf_4
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3984_ _3984_/A _4133_/A _3984_/C vssd1 vssd1 vccd1 vccd1 _3984_/X sky130_fd_sc_hd__and3_1
X_5723_ _5748_/A _5748_/B _5748_/C vssd1 vssd1 vccd1 vccd1 _5723_/Y sky130_fd_sc_hd__nand3_1
X_5654_ _5654_/A _6076_/A _5994_/B vssd1 vssd1 vccd1 vccd1 _5654_/X sky130_fd_sc_hd__and3_1
XFILLER_30_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4605_ _4605_/A _4605_/B _4605_/C vssd1 vssd1 vccd1 vccd1 _4606_/B sky130_fd_sc_hd__nand3_1
X_5585_ _5585_/A _5585_/B vssd1 vssd1 vccd1 vccd1 _5588_/A sky130_fd_sc_hd__nand2_2
X_4536_ _4531_/Y _4536_/B _4536_/C vssd1 vssd1 vccd1 vccd1 _4557_/B sky130_fd_sc_hd__nand3b_2
X_4467_ _4467_/A vssd1 vssd1 vccd1 vccd1 _4641_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6206_ _6244_/B _6206_/B _6206_/C vssd1 vssd1 vccd1 vccd1 _6208_/A sky130_fd_sc_hd__nand3_2
X_4398_ _4397_/C _4397_/A _4397_/B vssd1 vssd1 vccd1 vccd1 _4400_/B sky130_fd_sc_hd__a21o_1
X_3418_ _3418_/A _3866_/A vssd1 vssd1 vccd1 vccd1 _3419_/B sky130_fd_sc_hd__nand2_2
XFILLER_85_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6137_ _6137_/A _6137_/B _6137_/C _6137_/D vssd1 vssd1 vccd1 vccd1 _6138_/B sky130_fd_sc_hd__and4_2
X_3349_ _3287_/X _3345_/Y _3347_/Y _3440_/B vssd1 vssd1 vccd1 vccd1 _3349_/Y sky130_fd_sc_hd__o2bb2ai_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6068_ _6072_/A _6068_/B _6072_/B vssd1 vssd1 vccd1 vccd1 _6068_/X sky130_fd_sc_hd__and3_1
X_5019_ _5006_/Y _5007_/Y _5010_/X vssd1 vssd1 vccd1 vccd1 _5019_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5370_ _5603_/C _5046_/B _5239_/Y _5240_/X _5241_/X vssd1 vssd1 vccd1 vccd1 _5370_/X
+ sky130_fd_sc_hd__o221a_2
X_4321_ _4321_/A _4321_/B vssd1 vssd1 vccd1 vccd1 _4322_/C sky130_fd_sc_hd__nand2_1
X_4252_ _4252_/A vssd1 vssd1 vccd1 vccd1 _5286_/B sky130_fd_sc_hd__buf_2
X_3203_ _3170_/A _3170_/B _3201_/A _3201_/B _6297_/A vssd1 vssd1 vccd1 vccd1 _3245_/A
+ sky130_fd_sc_hd__o221ai_4
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4183_ _3791_/C _4179_/X _4197_/B _4182_/Y vssd1 vssd1 vccd1 vccd1 _4213_/A sky130_fd_sc_hd__a22o_1
X_3134_ _4067_/A vssd1 vssd1 vccd1 vccd1 _3218_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3967_ _4143_/A _4143_/B _3968_/A vssd1 vssd1 vccd1 vccd1 _4010_/A sky130_fd_sc_hd__o21a_1
XFILLER_23_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5706_ _5442_/C _5411_/C _5688_/A _5917_/A vssd1 vssd1 vccd1 vccd1 _5706_/Y sky130_fd_sc_hd__a22oi_2
X_3898_ _5066_/A _5068_/B _4931_/A _4229_/B vssd1 vssd1 vccd1 vccd1 _3898_/X sky130_fd_sc_hd__and4_2
X_5637_ _5640_/C _5640_/D _5638_/A vssd1 vssd1 vccd1 vccd1 _5639_/B sky130_fd_sc_hd__a21o_1
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5568_ _5568_/A vssd1 vssd1 vccd1 vccd1 _5625_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4519_ _4519_/A _4519_/B vssd1 vssd1 vccd1 vccd1 _4519_/X sky130_fd_sc_hd__and2_1
X_5499_ _5337_/X _5335_/B _5340_/Y vssd1 vssd1 vccd1 vccd1 _5499_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4870_ _4858_/Y _4866_/X _4867_/Y _4869_/X vssd1 vssd1 vccd1 vccd1 _4871_/A sky130_fd_sc_hd__o211ai_1
XFILLER_60_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3821_ _3782_/X _3817_/Y _3837_/B _3837_/A vssd1 vssd1 vccd1 vccd1 _3821_/X sky130_fd_sc_hd__o211a_1
XFILLER_32_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3752_ _3810_/A vssd1 vssd1 vccd1 vccd1 _3752_/X sky130_fd_sc_hd__buf_2
XFILLER_9_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3683_ _3667_/X _3685_/B _3684_/A _3684_/B vssd1 vssd1 vccd1 vccd1 _3699_/A sky130_fd_sc_hd__o2bb2ai_2
X_5422_ _5411_/X _5213_/X _5413_/A _5413_/B vssd1 vssd1 vccd1 vccd1 _5423_/D sky130_fd_sc_hd__o211ai_1
X_5353_ _5141_/C _6283_/C _5007_/A _5348_/X vssd1 vssd1 vccd1 vccd1 _5354_/C sky130_fd_sc_hd__a31o_1
X_4304_ _4308_/A _4308_/B _4303_/Y vssd1 vssd1 vccd1 vccd1 _4304_/X sky130_fd_sc_hd__a21o_1
X_5284_ _5285_/A _5541_/A _5284_/C _5284_/D vssd1 vssd1 vccd1 vccd1 _5296_/D sky130_fd_sc_hd__nand4_4
X_4235_ _5251_/A _4235_/B _5530_/A _5037_/B vssd1 vssd1 vccd1 vccd1 _4235_/Y sky130_fd_sc_hd__nand4_2
X_4166_ _4166_/A _4166_/B _4520_/A vssd1 vssd1 vccd1 vccd1 _4520_/B sky130_fd_sc_hd__nand3_1
XFILLER_28_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4097_ _4097_/A _4097_/B vssd1 vssd1 vccd1 vccd1 _4097_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4999_ _4990_/Y _4985_/Y _4979_/Y vssd1 vssd1 vccd1 vccd1 _5021_/C sky130_fd_sc_hd__a21o_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4020_ _4020_/A _4020_/B vssd1 vssd1 vccd1 vccd1 _4020_/Y sky130_fd_sc_hd__nand2_2
XFILLER_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5971_ _5971_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5984_/A sky130_fd_sc_hd__nand2_2
X_4922_ _4922_/A _5100_/A _5100_/B vssd1 vssd1 vccd1 vccd1 _4922_/X sky130_fd_sc_hd__and3_1
XFILLER_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4853_ _4853_/A _4853_/B vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__nand2_1
X_3804_ _3626_/X _3803_/X _3806_/A vssd1 vssd1 vccd1 vccd1 _3804_/X sky130_fd_sc_hd__o21a_1
X_4784_ _4784_/A _4784_/B _5436_/A _5582_/A vssd1 vssd1 vccd1 vccd1 _4786_/B sky130_fd_sc_hd__nand4_1
X_3735_ _3609_/X _3610_/Y _3733_/Y _3734_/X vssd1 vssd1 vccd1 vccd1 _3856_/B sky130_fd_sc_hd__a2bb2oi_2
X_5405_ _5407_/A _5407_/B _5656_/A _5407_/C vssd1 vssd1 vccd1 vccd1 _5405_/Y sky130_fd_sc_hd__nand4_4
X_3666_ _3666_/A _3666_/B _3666_/C vssd1 vssd1 vccd1 vccd1 _3685_/A sky130_fd_sc_hd__nand3_2
X_3597_ _3597_/A _3597_/B vssd1 vssd1 vccd1 vccd1 _3597_/Y sky130_fd_sc_hd__nand2_1
X_5336_ _5336_/A vssd1 vssd1 vccd1 vccd1 _5336_/Y sky130_fd_sc_hd__inv_2
X_5267_ _5420_/A _5267_/B vssd1 vssd1 vccd1 vccd1 _5424_/A sky130_fd_sc_hd__nand2_1
X_4218_ _4516_/C _4209_/B _4194_/Y _4198_/Y _4213_/Y vssd1 vssd1 vccd1 vccd1 _4220_/C
+ sky130_fd_sc_hd__o221ai_1
X_5198_ _5182_/B _5182_/C _5182_/A vssd1 vssd1 vccd1 vccd1 _5355_/A sky130_fd_sc_hd__a21boi_1
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4149_ _4142_/Y _4144_/X _4123_/Y _4125_/Y _4317_/A vssd1 vssd1 vccd1 vccd1 _4150_/C
+ sky130_fd_sc_hd__o221ai_1
XFILLER_28_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3520_ _5663_/A vssd1 vssd1 vccd1 vccd1 _5850_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3451_ _3342_/B _3530_/A _3204_/B _4422_/C _3443_/X vssd1 vssd1 vccd1 vccd1 _3452_/C
+ sky130_fd_sc_hd__o2111ai_2
X_6170_ _6170_/A _6170_/B _6170_/C _6170_/D vssd1 vssd1 vccd1 vccd1 _6198_/A sky130_fd_sc_hd__and4_1
X_3382_ _3382_/A vssd1 vssd1 vccd1 vccd1 _3484_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5121_ _5037_/B _4530_/C _5701_/A _5530_/A vssd1 vssd1 vccd1 vccd1 _5121_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_69_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5052_ _4868_/Y _5051_/Y _5087_/B vssd1 vssd1 vccd1 vccd1 _5082_/B sky130_fd_sc_hd__o21ai_1
X_4003_ _3998_/A _3998_/C _4163_/C _4163_/D vssd1 vssd1 vccd1 vccd1 _4004_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5954_ _5877_/X _5869_/Y _5900_/Y vssd1 vssd1 vccd1 vccd1 _5956_/A sky130_fd_sc_hd__o21a_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5885_ _5761_/A _5761_/B _5761_/C _5766_/C vssd1 vssd1 vccd1 vccd1 _5885_/Y sky130_fd_sc_hd__a31oi_2
X_4905_ _5401_/A _5449_/A _4903_/Y _4904_/Y vssd1 vssd1 vccd1 vccd1 _4913_/B sky130_fd_sc_hd__a22o_1
XFILLER_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4836_ _4671_/A _4671_/B _4671_/C _4679_/B _4680_/C vssd1 vssd1 vccd1 vccd1 _4839_/A
+ sky130_fd_sc_hd__a32oi_4
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4767_ _4599_/B _4606_/C _4577_/Y _4574_/Y vssd1 vssd1 vccd1 vccd1 _4772_/A sky130_fd_sc_hd__o2bb2ai_1
X_3718_ _3667_/X _3685_/B _3710_/X _3717_/X vssd1 vssd1 vccd1 vccd1 _3719_/C sky130_fd_sc_hd__o2bb2ai_1
X_4698_ _4698_/A _4928_/A vssd1 vssd1 vccd1 vccd1 _4698_/Y sky130_fd_sc_hd__nor2_4
XFILLER_20_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3649_ _4407_/A vssd1 vssd1 vccd1 vccd1 _5123_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5319_ _5366_/A _5366_/B vssd1 vssd1 vccd1 vccd1 _5328_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_9 _5780_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5670_ _5580_/Y _5832_/A _5994_/B _6077_/B _5852_/A vssd1 vssd1 vccd1 vccd1 _5671_/C
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4621_ _4621_/A _4621_/B _4621_/C _5401_/A vssd1 vssd1 vccd1 vccd1 _4623_/B sky130_fd_sc_hd__nand4_2
XFILLER_30_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4552_ _4531_/Y _4548_/X _4536_/C vssd1 vssd1 vccd1 vccd1 _4557_/A sky130_fd_sc_hd__o21bai_4
X_4483_ _4424_/X _4422_/X _4420_/X _4414_/X vssd1 vssd1 vccd1 vccd1 _4484_/B sky130_fd_sc_hd__o211ai_1
X_3503_ _3423_/Y _3502_/Y _3421_/Y vssd1 vssd1 vccd1 vccd1 _3509_/B sky130_fd_sc_hd__o21ai_2
X_6222_ _6222_/A _6222_/B vssd1 vssd1 vccd1 vccd1 _6224_/B sky130_fd_sc_hd__nor2_1
X_3434_ input7/X vssd1 vssd1 vccd1 vccd1 _4861_/A sky130_fd_sc_hd__buf_4
X_6153_ _6147_/Y _6150_/Y _6152_/Y vssd1 vssd1 vccd1 vccd1 _6153_/Y sky130_fd_sc_hd__o21ai_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _4956_/A _5374_/A vssd1 vssd1 vccd1 vccd1 _3368_/B sky130_fd_sc_hd__nand2_2
X_6084_ _6084_/A _6084_/B vssd1 vssd1 vccd1 vccd1 _6084_/Y sky130_fd_sc_hd__xnor2_1
X_5104_ _5104_/A vssd1 vssd1 vccd1 vccd1 _5203_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _4747_/A _3280_/X _3215_/B _3342_/A _3287_/X vssd1 vssd1 vccd1 vccd1 _3296_/Y
+ sky130_fd_sc_hd__o221ai_4
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5040_/A _5040_/B _5032_/B vssd1 vssd1 vccd1 vccd1 _5035_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5937_ _5937_/A vssd1 vssd1 vccd1 vccd1 _5942_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5868_ _5868_/A _5868_/B _5868_/C vssd1 vssd1 vccd1 vccd1 _5912_/A sky130_fd_sc_hd__and3_1
XFILLER_21_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5799_ _5799_/A _5799_/B vssd1 vssd1 vccd1 vccd1 _5799_/Y sky130_fd_sc_hd__nand2_1
X_4819_ _4819_/A _4819_/B _4819_/C vssd1 vssd1 vccd1 vccd1 _4819_/Y sky130_fd_sc_hd__nand3_4
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput57 _3171_/Y vssd1 vssd1 vccd1 vccd1 r[2] sky130_fd_sc_hd__buf_2
Xoutput46 _6297_/Y vssd1 vssd1 vccd1 vccd1 r[1] sky130_fd_sc_hd__buf_2
Xoutput35 _3150_/C vssd1 vssd1 vccd1 vccd1 r[0] sky130_fd_sc_hd__buf_2
Xoutput68 _3745_/X vssd1 vssd1 vccd1 vccd1 r[9] sky130_fd_sc_hd__buf_2
XFILLER_88_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3150_ _3190_/C _4832_/C _3150_/C vssd1 vssd1 vccd1 vccd1 _3151_/A sky130_fd_sc_hd__and3_1
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5722_ _5584_/A _5584_/B _5584_/C _5608_/C _5721_/X vssd1 vssd1 vccd1 vccd1 _5748_/C
+ sky130_fd_sc_hd__a32oi_4
X_3983_ _3882_/B _3882_/C _3980_/Y _4043_/C vssd1 vssd1 vccd1 vccd1 _3984_/A sky130_fd_sc_hd__o22ai_2
X_5653_ _5925_/B vssd1 vssd1 vccd1 vccd1 _6076_/A sky130_fd_sc_hd__clkbuf_2
X_5584_ _5584_/A _5584_/B _5584_/C vssd1 vssd1 vccd1 vccd1 _5608_/B sky130_fd_sc_hd__nand3_2
X_4604_ _4576_/B _4576_/C _4576_/A vssd1 vssd1 vccd1 vccd1 _4605_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4535_ _4366_/Y _4368_/Y _4363_/Y vssd1 vssd1 vccd1 vccd1 _4536_/C sky130_fd_sc_hd__o21ai_1
XFILLER_7_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4466_ _4466_/A _4466_/B _4466_/C vssd1 vssd1 vccd1 vccd1 _4467_/A sky130_fd_sc_hd__nand3_1
X_6205_ _6236_/C _6205_/B _6205_/C vssd1 vssd1 vccd1 vccd1 _6206_/C sky130_fd_sc_hd__and3_1
X_4397_ _4397_/A _4397_/B _4397_/C vssd1 vssd1 vccd1 vccd1 _4400_/A sky130_fd_sc_hd__nand3_2
X_3417_ _3772_/A vssd1 vssd1 vccd1 vccd1 _3418_/A sky130_fd_sc_hd__clkbuf_4
X_6136_ _6137_/C _4830_/A _6137_/D _6137_/A vssd1 vssd1 vccd1 vccd1 _6138_/A sky130_fd_sc_hd__a22oi_2
X_3348_ _3348_/A _3348_/B vssd1 vssd1 vccd1 vccd1 _3440_/B sky130_fd_sc_hd__nand2_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3279_ _4019_/A vssd1 vssd1 vccd1 vccd1 _3280_/A sky130_fd_sc_hd__inv_2
X_6067_ _6072_/A _6072_/B _6068_/B vssd1 vssd1 vccd1 vccd1 _6067_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_85_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5018_ _5018_/A vssd1 vssd1 vccd1 vccd1 _5018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4320_ _4226_/B _4225_/A _4313_/A vssd1 vssd1 vccd1 vccd1 _4321_/A sky130_fd_sc_hd__a21o_1
XFILLER_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4251_ _5245_/A _5068_/B _5123_/A _4777_/D vssd1 vssd1 vccd1 vccd1 _4251_/Y sky130_fd_sc_hd__nand4_2
XFILLER_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3202_ _3202_/A _3202_/B vssd1 vssd1 vccd1 vccd1 _3202_/Y sky130_fd_sc_hd__xnor2_4
X_4182_ _4182_/A _4182_/B vssd1 vssd1 vccd1 vccd1 _4182_/Y sky130_fd_sc_hd__nand2_2
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3133_ _5045_/A vssd1 vssd1 vccd1 vccd1 _4067_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3966_ _3966_/A _3966_/B _6127_/A _6165_/A vssd1 vssd1 vccd1 vccd1 _3968_/A sky130_fd_sc_hd__nand4_4
XFILLER_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5705_ _5697_/A _5697_/B _5704_/Y vssd1 vssd1 vccd1 vccd1 _5799_/B sky130_fd_sc_hd__o21ai_1
XFILLER_10_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5636_ _5640_/A _5640_/B vssd1 vssd1 vccd1 vccd1 _5638_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3897_ _3897_/A vssd1 vssd1 vccd1 vccd1 _5068_/B sky130_fd_sc_hd__clkbuf_4
X_5567_ _5567_/A _5567_/B _5567_/C vssd1 vssd1 vccd1 vccd1 _5568_/A sky130_fd_sc_hd__nand3_1
X_5498_ _5327_/Y _5495_/Y _5502_/A _5525_/A vssd1 vssd1 vccd1 vccd1 _5498_/X sky130_fd_sc_hd__o211a_1
X_4518_ _4842_/A _4842_/B vssd1 vssd1 vccd1 vccd1 _4518_/X sky130_fd_sc_hd__and2_1
X_4449_ _5065_/A _5206_/A vssd1 vssd1 vccd1 vccd1 _4449_/Y sky130_fd_sc_hd__nand2_1
X_6119_ _6108_/A _6108_/B _6108_/C vssd1 vssd1 vccd1 vccd1 _6119_/Y sky130_fd_sc_hd__a21oi_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3820_ _3822_/C _3822_/B _3808_/A _3808_/B vssd1 vssd1 vccd1 vccd1 _3837_/A sky130_fd_sc_hd__o2bb2ai_2
X_3751_ _3755_/A _3755_/B _3755_/C vssd1 vssd1 vccd1 vccd1 _3810_/A sky130_fd_sc_hd__a21oi_1
X_3682_ _3611_/X _3679_/Y _3681_/X _3676_/Y vssd1 vssd1 vccd1 vccd1 _3684_/B sky130_fd_sc_hd__o211a_1
X_5421_ _5414_/Y _5415_/X _5413_/C vssd1 vssd1 vccd1 vccd1 _5423_/C sky130_fd_sc_hd__o21ai_1
X_5352_ _5352_/A vssd1 vssd1 vccd1 vccd1 _6283_/C sky130_fd_sc_hd__clkbuf_4
X_4303_ _4308_/C _4308_/D vssd1 vssd1 vccd1 vccd1 _4303_/Y sky130_fd_sc_hd__nand2_1
X_5283_ _5485_/A _5485_/B _5484_/A vssd1 vssd1 vccd1 vccd1 _5283_/Y sky130_fd_sc_hd__nand3_2
XFILLER_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4234_ _4234_/A vssd1 vssd1 vccd1 vccd1 _5037_/B sky130_fd_sc_hd__clkbuf_4
X_4165_ _4165_/A vssd1 vssd1 vccd1 vccd1 _4520_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4096_ _4096_/A _4097_/A _4097_/B vssd1 vssd1 vccd1 vccd1 _4096_/X sky130_fd_sc_hd__and3_1
XFILLER_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4998_ _4927_/Y _4973_/Y _4979_/Y _4985_/Y vssd1 vssd1 vccd1 vccd1 _5021_/B sky130_fd_sc_hd__o211ai_4
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3949_ _4936_/B vssd1 vssd1 vccd1 vccd1 _5704_/B sky130_fd_sc_hd__buf_2
X_5619_ _5430_/A _5614_/Y _5611_/A _5611_/B vssd1 vssd1 vccd1 vccd1 _5619_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_58_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ _6058_/A _5969_/B _5969_/C vssd1 vssd1 vccd1 vccd1 _5971_/B sky130_fd_sc_hd__a21o_1
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4921_ _4921_/A _4981_/A vssd1 vssd1 vccd1 vccd1 _4972_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4852_ _4852_/A _5230_/A vssd1 vssd1 vccd1 vccd1 _4853_/B sky130_fd_sc_hd__nand2_2
X_3803_ _3803_/A _3803_/B _5831_/A _5669_/A vssd1 vssd1 vccd1 vccd1 _3803_/X sky130_fd_sc_hd__and4_1
XFILLER_20_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4783_ _4935_/A vssd1 vssd1 vccd1 vccd1 _5436_/A sky130_fd_sc_hd__buf_2
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3734_ _3835_/A _3836_/A _3835_/B vssd1 vssd1 vccd1 vccd1 _3734_/X sky130_fd_sc_hd__a21o_1
X_3665_ _3441_/X _3669_/A _3530_/B _3747_/A _3761_/A vssd1 vssd1 vccd1 vccd1 _3666_/C
+ sky130_fd_sc_hd__o221ai_1
X_5404_ _5580_/A _5404_/B _5794_/C _5918_/B vssd1 vssd1 vccd1 vccd1 _5407_/B sky130_fd_sc_hd__nand4_2
X_3596_ _3596_/A _3596_/B vssd1 vssd1 vccd1 vccd1 _3857_/B sky130_fd_sc_hd__nand2_2
XFILLER_87_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5335_ _5335_/A _5335_/B vssd1 vssd1 vccd1 vccd1 _5339_/B sky130_fd_sc_hd__nand2_1
X_5266_ _5420_/B _5420_/C vssd1 vssd1 vccd1 vccd1 _5267_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4217_ _4226_/B vssd1 vssd1 vccd1 vccd1 _4313_/B sky130_fd_sc_hd__clkbuf_1
X_5197_ _5197_/A vssd1 vssd1 vccd1 vccd1 _5197_/X sky130_fd_sc_hd__clkbuf_1
X_4148_ _4011_/X _3973_/B _3984_/X _3985_/Y vssd1 vssd1 vccd1 vccd1 _4150_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4079_ _4855_/B _5029_/B vssd1 vssd1 vccd1 vccd1 _4079_/Y sky130_fd_sc_hd__nand2_2
XFILLER_70_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3450_ _4363_/B vssd1 vssd1 vccd1 vccd1 _4422_/C sky130_fd_sc_hd__buf_4
X_3381_ _3398_/B _3381_/B _3381_/C vssd1 vssd1 vccd1 vccd1 _3382_/A sky130_fd_sc_hd__nand3b_1
XFILLER_69_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5120_ _5120_/A _5128_/B vssd1 vssd1 vccd1 vccd1 _5120_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5051_ _4734_/B _5059_/A _5237_/A _4432_/A vssd1 vssd1 vccd1 vccd1 _5051_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_84_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4002_ _4161_/A _4002_/B _4161_/B vssd1 vssd1 vccd1 vccd1 _4163_/D sky130_fd_sc_hd__nand3_1
XFILLER_84_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5953_ _5960_/A _5960_/B _5960_/C vssd1 vssd1 vccd1 vccd1 _5957_/C sky130_fd_sc_hd__nand3_1
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5884_ _5884_/A vssd1 vssd1 vccd1 vccd1 _5884_/Y sky130_fd_sc_hd__inv_2
X_4904_ _5209_/A _4904_/B _5223_/A _5448_/B vssd1 vssd1 vccd1 vccd1 _4904_/Y sky130_fd_sc_hd__nand4_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4835_ _5190_/A _5190_/B _4834_/X vssd1 vssd1 vccd1 vccd1 _4845_/A sky130_fd_sc_hd__o21ai_1
X_4766_ _4766_/A vssd1 vssd1 vccd1 vccd1 _4801_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3717_ _3713_/Y _3714_/X _5007_/A _5858_/C vssd1 vssd1 vccd1 vccd1 _3717_/X sky130_fd_sc_hd__o211a_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4697_ _4935_/B _4935_/C vssd1 vssd1 vccd1 vccd1 _4928_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3648_ _4852_/A vssd1 vssd1 vccd1 vccd1 _5048_/A sky130_fd_sc_hd__buf_4
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3579_ _3574_/X _3575_/Y _3609_/B _3609_/C vssd1 vssd1 vccd1 vccd1 _3607_/C sky130_fd_sc_hd__o211ai_4
X_5318_ _5277_/Y _5283_/Y _5316_/Y _5317_/X vssd1 vssd1 vccd1 vccd1 _5323_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5249_ _5250_/A _5246_/X _5248_/Y vssd1 vssd1 vccd1 vccd1 _5249_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _5435_/A _5582_/A _4621_/A _4621_/B vssd1 vssd1 vccd1 vccd1 _4623_/A sky130_fd_sc_hd__a22o_1
X_4551_ _4414_/X _4550_/X _4420_/X vssd1 vssd1 vccd1 vccd1 _4551_/Y sky130_fd_sc_hd__a21boi_4
X_4482_ _4422_/A _4231_/Y _4414_/A _4420_/A vssd1 vssd1 vccd1 vccd1 _4484_/A sky130_fd_sc_hd__a22o_1
X_3502_ _5597_/A _5134_/A _5596_/B _3803_/B vssd1 vssd1 vccd1 vccd1 _3502_/Y sky130_fd_sc_hd__a22oi_2
X_6221_ _5981_/A _5981_/B _6220_/Y vssd1 vssd1 vccd1 vccd1 _6221_/Y sky130_fd_sc_hd__a21oi_2
X_3433_ _4571_/A _4935_/B vssd1 vssd1 vccd1 vccd1 _3433_/Y sky130_fd_sc_hd__nand2_1
X_6152_ _6147_/Y _6151_/Y _6149_/Y vssd1 vssd1 vccd1 vccd1 _6152_/Y sky130_fd_sc_hd__o21bai_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5102_/Y _4981_/B _4981_/C vssd1 vssd1 vccd1 vccd1 _5103_/Y sky130_fd_sc_hd__a21boi_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _4019_/A vssd1 vssd1 vccd1 vccd1 _4956_/A sky130_fd_sc_hd__clkbuf_2
X_6083_ _6089_/C _6089_/B _6087_/A _6087_/B vssd1 vssd1 vccd1 vccd1 _6083_/Y sky130_fd_sc_hd__nand4_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _3295_/A _3295_/B _3295_/C vssd1 vssd1 vccd1 vccd1 _3300_/C sky130_fd_sc_hd__nand3_2
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5034_/A _5034_/B vssd1 vssd1 vccd1 vccd1 _5040_/B sky130_fd_sc_hd__nor2_1
XFILLER_65_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5936_ _5936_/A _5942_/A vssd1 vssd1 vccd1 vccd1 _5940_/A sky130_fd_sc_hd__nand2_1
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5867_ _5867_/A _6236_/B vssd1 vssd1 vccd1 vccd1 _5868_/C sky130_fd_sc_hd__nor2_1
X_5798_ _5793_/A _5793_/B _5789_/Y vssd1 vssd1 vccd1 vccd1 _5798_/Y sky130_fd_sc_hd__o21ai_1
X_4818_ _4817_/A _4817_/B _4822_/B _4816_/A vssd1 vssd1 vccd1 vccd1 _4819_/C sky130_fd_sc_hd__a22o_1
XFILLER_31_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4749_ _4579_/Y _4743_/X _4745_/Y _4748_/Y vssd1 vssd1 vccd1 vccd1 _4749_/Y sky130_fd_sc_hd__o211ai_2
Xoutput58 _6251_/Y vssd1 vssd1 vccd1 vccd1 r[30] sky130_fd_sc_hd__buf_2
Xoutput47 _5523_/X vssd1 vssd1 vccd1 vccd1 r[20] sky130_fd_sc_hd__buf_2
Xoutput36 _3859_/X vssd1 vssd1 vccd1 vccd1 r[10] sky130_fd_sc_hd__buf_2
XFILLER_88_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3982_ _3882_/C _3981_/Y _3882_/B vssd1 vssd1 vccd1 vccd1 _4043_/C sky130_fd_sc_hd__o21ai_4
XFILLER_35_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5721_ _5208_/B _5399_/Y _5405_/Y vssd1 vssd1 vccd1 vccd1 _5721_/X sky130_fd_sc_hd__o21a_1
XFILLER_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5652_ _5850_/A _5833_/B _6077_/B _6071_/A vssd1 vssd1 vccd1 vccd1 _5652_/X sky130_fd_sc_hd__and4_1
X_5583_ _5585_/B _5583_/B vssd1 vssd1 vccd1 vccd1 _5584_/C sky130_fd_sc_hd__nand2_1
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4603_ _4267_/Y _4568_/A _4443_/Y _4575_/Y vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__o22a_1
X_4534_ _4365_/B _4533_/X _4939_/A _4038_/B _4529_/Y vssd1 vssd1 vccd1 vccd1 _4536_/B
+ sky130_fd_sc_hd__o2111ai_1
X_4465_ _4464_/X _4266_/Y _4270_/Y _4294_/B _4294_/C vssd1 vssd1 vccd1 vccd1 _4466_/C
+ sky130_fd_sc_hd__a32oi_4
X_6204_ _6203_/X _6202_/A _5352_/A _6072_/C vssd1 vssd1 vccd1 vccd1 _6206_/B sky130_fd_sc_hd__a2bb2o_1
X_4396_ _4399_/A _4399_/B _4394_/X _4395_/Y vssd1 vssd1 vccd1 vccd1 _4495_/A sky130_fd_sc_hd__o22ai_4
X_3416_ _4956_/A _4454_/B vssd1 vssd1 vccd1 vccd1 _3419_/A sky130_fd_sc_hd__nand2_1
X_6135_ _6170_/B _6134_/C _6170_/C _6170_/A vssd1 vssd1 vccd1 vccd1 _6137_/A sky130_fd_sc_hd__a22o_1
X_3347_ _3270_/B _4958_/B _5299_/A _3458_/A vssd1 vssd1 vccd1 vccd1 _3347_/Y sky130_fd_sc_hd__a22oi_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _6165_/B _6071_/A vssd1 vssd1 vccd1 vccd1 _6068_/B sky130_fd_sc_hd__and2_1
X_5017_ _5017_/A _5017_/B vssd1 vssd1 vccd1 vccd1 _5018_/A sky130_fd_sc_hd__and2_2
X_3278_ _3894_/A vssd1 vssd1 vccd1 vccd1 _4747_/A sky130_fd_sc_hd__buf_4
XFILLER_26_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5919_ _5919_/A _5919_/B vssd1 vssd1 vccd1 vccd1 _5920_/B sky130_fd_sc_hd__nand2_1
XFILLER_42_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _4302_/C _4302_/D _4250_/C vssd1 vssd1 vccd1 vccd1 _4250_/X sky130_fd_sc_hd__and3_1
X_4181_ _4184_/A _5696_/A vssd1 vssd1 vccd1 vccd1 _4182_/B sky130_fd_sc_hd__nand2_2
X_3201_ _3201_/A _3201_/B vssd1 vssd1 vccd1 vccd1 _3202_/B sky130_fd_sc_hd__or2_2
X_3132_ input1/X vssd1 vssd1 vccd1 vccd1 _5045_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3965_ _5919_/A vssd1 vssd1 vccd1 vccd1 _6127_/A sky130_fd_sc_hd__buf_2
X_5704_ _5704_/A _5704_/B vssd1 vssd1 vccd1 vccd1 _5704_/Y sky130_fd_sc_hd__nand2_1
X_3896_ _4096_/A _4097_/A _4097_/B vssd1 vssd1 vccd1 vccd1 _3927_/A sky130_fd_sc_hd__nand3_1
X_5635_ _5635_/A _5635_/B _5635_/C vssd1 vssd1 vccd1 vccd1 _5640_/D sky130_fd_sc_hd__nand3_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5566_ _5566_/A vssd1 vssd1 vccd1 vccd1 _5625_/A sky130_fd_sc_hd__clkbuf_2
X_5497_ _5502_/A _5525_/A _5502_/C vssd1 vssd1 vccd1 vccd1 _5497_/Y sky130_fd_sc_hd__a21oi_1
X_4517_ _4519_/B _4517_/B _4517_/C vssd1 vssd1 vccd1 vccd1 _4842_/B sky130_fd_sc_hd__nand3b_2
X_4448_ _4874_/A _4901_/B vssd1 vssd1 vccd1 vccd1 _4592_/A sky130_fd_sc_hd__nand2_1
X_4379_ _4359_/X _4362_/X _4378_/Y vssd1 vssd1 vccd1 vccd1 _4397_/A sky130_fd_sc_hd__o21ai_2
X_6118_ _6118_/A _6118_/B vssd1 vssd1 vccd1 vccd1 _6118_/X sky130_fd_sc_hd__xor2_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _6049_/A _6049_/B vssd1 vssd1 vccd1 vccd1 _6051_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3750_ _4744_/A _4930_/A vssd1 vssd1 vccd1 vccd1 _3755_/C sky130_fd_sc_hd__and2_1
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3681_ _4184_/A _4880_/A vssd1 vssd1 vccd1 vccd1 _3681_/X sky130_fd_sc_hd__and2_1
X_5420_ _5420_/A _5420_/B _5420_/C vssd1 vssd1 vccd1 vccd1 _5420_/X sky130_fd_sc_hd__and3_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5351_ _5351_/A vssd1 vssd1 vccd1 vccd1 _5513_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5282_ _5427_/A _5427_/B _5490_/A _5431_/A vssd1 vssd1 vccd1 vccd1 _5484_/A sky130_fd_sc_hd__nand4_2
X_4302_ _4302_/A _4302_/B _4302_/C _4302_/D vssd1 vssd1 vccd1 vccd1 _4308_/D sky130_fd_sc_hd__nand4_2
X_4233_ _5119_/A vssd1 vssd1 vccd1 vccd1 _5530_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4164_ _4163_/B _3998_/D _4163_/Y _3859_/B vssd1 vssd1 vccd1 vccd1 _4164_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_95_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4095_ _4095_/A _4095_/B _4095_/C vssd1 vssd1 vccd1 vccd1 _4124_/C sky130_fd_sc_hd__nand3_4
XFILLER_67_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4997_ _4822_/A _4822_/C _4995_/Y _4996_/Y vssd1 vssd1 vccd1 vccd1 _5020_/B sky130_fd_sc_hd__o2bb2ai_4
XFILLER_23_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3948_ input3/X vssd1 vssd1 vccd1 vccd1 _4936_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3879_ _5134_/A _5831_/A _5669_/A _3555_/A vssd1 vssd1 vccd1 vccd1 _3879_/Y sky130_fd_sc_hd__a22oi_1
X_5618_ _5618_/A _5625_/C _5625_/D vssd1 vssd1 vccd1 vccd1 _5622_/B sky130_fd_sc_hd__nand3_1
X_5549_ _5549_/A _5549_/B _5549_/C vssd1 vssd1 vccd1 vccd1 _5694_/C sky130_fd_sc_hd__nand3_1
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4920_ _4912_/Y _4922_/A _4919_/Y vssd1 vssd1 vccd1 vccd1 _4981_/A sky130_fd_sc_hd__a21oi_1
XFILLER_52_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4851_ _4819_/Y _4850_/X _4824_/Y vssd1 vssd1 vccd1 vccd1 _5012_/A sky130_fd_sc_hd__a21boi_2
X_3802_ _5575_/A vssd1 vssd1 vccd1 vccd1 _5669_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4782_ _5532_/A _4110_/B _4784_/A _4784_/B vssd1 vssd1 vccd1 vccd1 _4786_/A sky130_fd_sc_hd__a22o_1
X_3733_ _3835_/A _3836_/A _3835_/B vssd1 vssd1 vccd1 vccd1 _3733_/Y sky130_fd_sc_hd__nand3_2
X_3664_ _4855_/B _4930_/A _4234_/A _4855_/A vssd1 vssd1 vccd1 vccd1 _3761_/A sky130_fd_sc_hd__a22o_2
X_5403_ _5403_/A _5403_/B vssd1 vssd1 vccd1 vccd1 _5407_/A sky130_fd_sc_hd__nand2_1
X_3595_ _3596_/A _3596_/B _3597_/A vssd1 vssd1 vccd1 vccd1 _6294_/B sky130_fd_sc_hd__a21o_1
X_5334_ _5336_/A _5163_/C _5333_/X vssd1 vssd1 vccd1 vccd1 _5335_/B sky130_fd_sc_hd__a21o_1
X_5265_ _5594_/A _5917_/C _5263_/A _5263_/B vssd1 vssd1 vccd1 vccd1 _5420_/C sky130_fd_sc_hd__a22o_2
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5196_ _5196_/A _5196_/B vssd1 vssd1 vccd1 vccd1 _5197_/A sky130_fd_sc_hd__or2_4
X_4216_ _4399_/A _4210_/Y _4212_/Y _4215_/Y vssd1 vssd1 vccd1 vccd1 _4226_/B sky130_fd_sc_hd__o211ai_2
XFILLER_68_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4147_ _4317_/A _4141_/Y _4053_/Y _4054_/X vssd1 vssd1 vccd1 vccd1 _4150_/A sky130_fd_sc_hd__o2bb2ai_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4078_ _4078_/A vssd1 vssd1 vccd1 vccd1 _5029_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3380_ _3344_/Y _3349_/Y _3372_/B _3477_/A vssd1 vssd1 vccd1 vccd1 _3381_/C sky130_fd_sc_hd__o211ai_1
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5050_ _5081_/A _5081_/B _3189_/A _5599_/A vssd1 vssd1 vccd1 vccd1 _5082_/A sky130_fd_sc_hd__o2bb2ai_2
X_4001_ _4160_/A _4160_/B _4160_/C vssd1 vssd1 vccd1 vccd1 _4161_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5952_ _5952_/A _5952_/B _5952_/C vssd1 vssd1 vccd1 vccd1 _5960_/C sky130_fd_sc_hd__nand3_1
XFILLER_80_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4903_ _4903_/A _4903_/B vssd1 vssd1 vccd1 vccd1 _4903_/Y sky130_fd_sc_hd__nand2_2
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5883_ _5883_/A _5883_/B _5883_/C vssd1 vssd1 vccd1 vccd1 _5892_/B sky130_fd_sc_hd__nand3_1
XFILLER_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4834_ _4671_/A _4671_/B _4671_/C _4679_/B _4680_/C vssd1 vssd1 vccd1 vccd1 _4834_/X
+ sky130_fd_sc_hd__a32o_2
X_4765_ _4765_/A _4765_/B _4765_/C vssd1 vssd1 vccd1 vccd1 _4766_/A sky130_fd_sc_hd__nand3_1
X_3716_ _5263_/C vssd1 vssd1 vccd1 vccd1 _5858_/C sky130_fd_sc_hd__buf_4
X_4696_ _4423_/A _4935_/C _5448_/A _4532_/A vssd1 vssd1 vccd1 vccd1 _4703_/A sky130_fd_sc_hd__a22oi_2
X_3647_ input1/X vssd1 vssd1 vccd1 vccd1 _4852_/A sky130_fd_sc_hd__clkbuf_4
X_3578_ _3577_/B _3703_/B _3703_/A vssd1 vssd1 vccd1 vccd1 _3609_/C sky130_fd_sc_hd__a21o_2
XFILLER_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5317_ _5317_/A _5321_/B _5321_/C vssd1 vssd1 vccd1 vccd1 _5317_/X sky130_fd_sc_hd__and3_1
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6297_ _6297_/A _6297_/B vssd1 vssd1 vccd1 vccd1 _6297_/Y sky130_fd_sc_hd__nor2_4
XFILLER_75_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5248_ _5248_/A _5918_/B vssd1 vssd1 vccd1 vccd1 _5248_/Y sky130_fd_sc_hd__nand2_2
X_5179_ _5177_/Y _5178_/Y _5170_/B _5171_/C vssd1 vssd1 vccd1 vccd1 _5180_/C sky130_fd_sc_hd__o211ai_2
XFILLER_28_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4550_ _5511_/C _4422_/A _4422_/B _4424_/X vssd1 vssd1 vccd1 vccd1 _4550_/X sky130_fd_sc_hd__a31o_1
X_4481_ _4481_/A vssd1 vssd1 vccd1 vccd1 _4648_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3501_ _4956_/A vssd1 vssd1 vccd1 vccd1 _3803_/B sky130_fd_sc_hd__buf_4
X_6220_ _6220_/A _6220_/B vssd1 vssd1 vccd1 vccd1 _6220_/Y sky130_fd_sc_hd__nand2_1
X_3432_ _3774_/B vssd1 vssd1 vccd1 vccd1 _4935_/B sky130_fd_sc_hd__buf_2
X_6151_ _6151_/A _6151_/B vssd1 vssd1 vccd1 vccd1 _6151_/Y sky130_fd_sc_hd__nor2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _4540_/A _4235_/B vssd1 vssd1 vccd1 vccd1 _3368_/A sky130_fd_sc_hd__nand2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5099_/Y _5100_/Y _5101_/X vssd1 vssd1 vccd1 vccd1 _5102_/Y sky130_fd_sc_hd__o21ai_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6082_ _6079_/A _4830_/A _6084_/B vssd1 vssd1 vccd1 vccd1 _6087_/B sky130_fd_sc_hd__a21o_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _3223_/Y _3293_/Y _3229_/B vssd1 vssd1 vccd1 vccd1 _3295_/C sky130_fd_sc_hd__o21ai_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _4907_/X _5025_/B _5208_/A _4902_/A vssd1 vssd1 vccd1 vccd1 _5040_/A sky130_fd_sc_hd__o2bb2ai_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5935_ _5935_/A _5935_/B vssd1 vssd1 vccd1 vccd1 _5942_/A sky130_fd_sc_hd__nor2_2
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5866_ _5957_/A _5865_/B _5865_/C vssd1 vssd1 vccd1 vccd1 _5866_/Y sky130_fd_sc_hd__a21oi_1
X_4817_ _4817_/A _4817_/B _4822_/B _4822_/C vssd1 vssd1 vccd1 vccd1 _4819_/B sky130_fd_sc_hd__nand4_1
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5797_ _5823_/A vssd1 vssd1 vccd1 vccd1 _5816_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4748_ _4748_/A _4748_/B vssd1 vssd1 vccd1 vccd1 _4748_/Y sky130_fd_sc_hd__nand2_1
X_4679_ _4679_/A _4679_/B vssd1 vssd1 vccd1 vccd1 _4683_/A sky130_fd_sc_hd__nand2_1
Xoutput48 _5646_/Y vssd1 vssd1 vccd1 vccd1 r[21] sky130_fd_sc_hd__buf_2
Xoutput37 _4005_/Y vssd1 vssd1 vccd1 vccd1 r[11] sky130_fd_sc_hd__buf_2
Xoutput59 _6273_/Y vssd1 vssd1 vccd1 vccd1 r[31] sky130_fd_sc_hd__buf_2
XFILLER_88_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3981_ _3878_/A _3878_/B _3878_/C vssd1 vssd1 vccd1 vccd1 _3981_/Y sky130_fd_sc_hd__a21oi_2
X_5720_ _5724_/A _5728_/B _5733_/A _5733_/B vssd1 vssd1 vccd1 vccd1 _5748_/B sky130_fd_sc_hd__nand4_1
XFILLER_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5651_ _6002_/B vssd1 vssd1 vccd1 vccd1 _6071_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5582_ _5582_/A _5794_/C vssd1 vssd1 vccd1 vccd1 _5583_/B sky130_fd_sc_hd__and2_2
X_4602_ _4463_/B _4463_/C _4600_/X _4601_/Y vssd1 vssd1 vccd1 vccd1 _4607_/B sky130_fd_sc_hd__o2bb2ai_2
X_4533_ _4698_/A vssd1 vssd1 vccd1 vccd1 _4533_/X sky130_fd_sc_hd__clkbuf_2
X_6203_ _6203_/A _6233_/B _6203_/C _6203_/D vssd1 vssd1 vccd1 vccd1 _6203_/X sky130_fd_sc_hd__and4_1
X_4464_ _4064_/X _4079_/Y _4059_/Y _4063_/Y vssd1 vssd1 vccd1 vccd1 _4464_/X sky130_fd_sc_hd__o22a_1
X_4395_ _4397_/C _4397_/A _4397_/B vssd1 vssd1 vccd1 vccd1 _4395_/Y sky130_fd_sc_hd__a21oi_2
X_3415_ _4873_/A vssd1 vssd1 vccd1 vccd1 _4454_/B sky130_fd_sc_hd__buf_2
X_6134_ _6203_/A _6170_/B _6134_/C _6170_/C vssd1 vssd1 vccd1 vccd1 _6137_/D sky130_fd_sc_hd__nand4_1
X_3346_ _3542_/A vssd1 vssd1 vccd1 vccd1 _5299_/A sky130_fd_sc_hd__buf_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _6127_/A _6127_/B _6065_/C _6065_/D vssd1 vssd1 vccd1 vccd1 _6072_/B sky130_fd_sc_hd__nand4_2
XFILLER_85_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5016_ _5518_/A _4847_/B _5518_/B _4845_/B vssd1 vssd1 vccd1 vccd1 _5017_/B sky130_fd_sc_hd__o211ai_1
X_3277_ _3441_/A vssd1 vssd1 vccd1 vccd1 _3894_/A sky130_fd_sc_hd__clkbuf_4
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5918_ _6009_/A _5918_/B vssd1 vssd1 vccd1 vccd1 _5920_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5849_ _5659_/Y _5830_/X _5840_/Y _5848_/Y vssd1 vssd1 vccd1 vccd1 _5849_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_21_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4180_ _4366_/A _4958_/A _5792_/A _4363_/D vssd1 vssd1 vccd1 vccd1 _4197_/B sky130_fd_sc_hd__nand4_4
X_3200_ _3199_/A _3199_/B _3199_/C vssd1 vssd1 vccd1 vccd1 _3201_/B sky130_fd_sc_hd__a21oi_1
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3964_ _3964_/A _3964_/B _4362_/C _6010_/A vssd1 vssd1 vccd1 vccd1 _4143_/B sky130_fd_sc_hd__and4_2
X_5703_ _5703_/A _5703_/B _5703_/C vssd1 vssd1 vccd1 vccd1 _5724_/A sky130_fd_sc_hd__nand3_2
X_3895_ _3895_/A _3895_/B vssd1 vssd1 vccd1 vccd1 _4097_/B sky130_fd_sc_hd__nand2_2
X_5634_ _5634_/A _5634_/B _5634_/C _5634_/D vssd1 vssd1 vccd1 vccd1 _5635_/C sky130_fd_sc_hd__nand4_1
XFILLER_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5565_ _5567_/A _5567_/B _5567_/C vssd1 vssd1 vccd1 vccd1 _5566_/A sky130_fd_sc_hd__a21o_1
X_5496_ _5313_/A _5313_/B _5313_/C _5495_/Y vssd1 vssd1 vccd1 vccd1 _5502_/C sky130_fd_sc_hd__a31o_1
X_4516_ _4516_/A _4516_/B _4516_/C vssd1 vssd1 vccd1 vccd1 _4517_/C sky130_fd_sc_hd__nand3_1
X_4447_ _4460_/B vssd1 vssd1 vccd1 vccd1 _5453_/A sky130_fd_sc_hd__clkbuf_4
X_6117_ _5982_/B _6220_/A _6116_/X vssd1 vssd1 vccd1 vccd1 _6118_/B sky130_fd_sc_hd__a21boi_4
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4378_ _4367_/Y _4371_/Y _4377_/Y vssd1 vssd1 vccd1 vccd1 _4378_/Y sky130_fd_sc_hd__o21ai_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3329_ _4874_/A vssd1 vssd1 vccd1 vccd1 _5374_/A sky130_fd_sc_hd__clkbuf_4
X_6048_ _6048_/A _6048_/B vssd1 vssd1 vccd1 vccd1 _6049_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3680_ _4884_/A vssd1 vssd1 vccd1 vccd1 _4880_/A sky130_fd_sc_hd__clkbuf_4
X_5350_ _5350_/A _5364_/B vssd1 vssd1 vccd1 vccd1 _5355_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5281_ _5281_/A _5281_/B _5281_/C vssd1 vssd1 vccd1 vccd1 _5427_/B sky130_fd_sc_hd__nand3_2
X_4301_ _4302_/C _4302_/D _4250_/C vssd1 vssd1 vccd1 vccd1 _4308_/C sky130_fd_sc_hd__a21o_1
X_4232_ _5580_/A _4625_/A _5404_/B _5132_/B vssd1 vssd1 vccd1 vccd1 _4232_/Y sky130_fd_sc_hd__a22oi_4
X_4163_ _4163_/A _4163_/B _4163_/C _4163_/D vssd1 vssd1 vccd1 vccd1 _4163_/Y sky130_fd_sc_hd__nand4_2
XFILLER_95_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4094_ _4096_/A _4097_/A _4097_/B _4128_/A _4128_/B vssd1 vssd1 vccd1 vccd1 _4095_/C
+ sky130_fd_sc_hd__a32oi_4
XFILLER_67_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4996_ _4996_/A _4996_/B vssd1 vssd1 vccd1 vccd1 _4996_/Y sky130_fd_sc_hd__nand2_1
X_3947_ _4008_/A _4008_/B _4008_/C vssd1 vssd1 vccd1 vccd1 _3973_/B sky130_fd_sc_hd__nand3_2
X_3878_ _3878_/A _3878_/B _3878_/C vssd1 vssd1 vccd1 vccd1 _3882_/B sky130_fd_sc_hd__nand3_2
X_5617_ _5612_/X _5613_/Y _5614_/Y _5611_/A _5611_/B vssd1 vssd1 vccd1 vccd1 _5625_/D
+ sky130_fd_sc_hd__o2111ai_4
X_5548_ _5546_/Y _5547_/Y _5442_/Y vssd1 vssd1 vccd1 vccd1 _5549_/C sky130_fd_sc_hd__o21ai_2
X_5479_ _5479_/A _5479_/B vssd1 vssd1 vccd1 vccd1 _5634_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4850_ _4832_/A _6255_/B _4832_/C _4827_/X vssd1 vssd1 vccd1 vccd1 _4850_/X sky130_fd_sc_hd__a31o_1
X_3801_ _5029_/A vssd1 vssd1 vccd1 vccd1 _5575_/A sky130_fd_sc_hd__clkbuf_4
X_4781_ _4781_/A _4781_/B _4781_/C vssd1 vssd1 vccd1 vccd1 _4950_/A sky130_fd_sc_hd__nand3_4
X_3732_ _3732_/A _3845_/B vssd1 vssd1 vccd1 vccd1 _3835_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3663_ input1/X vssd1 vssd1 vccd1 vccd1 _4855_/A sky130_fd_sc_hd__buf_2
X_5402_ _5402_/A _5402_/B vssd1 vssd1 vccd1 vccd1 _5402_/Y sky130_fd_sc_hd__nand2_2
X_5333_ _5099_/Y _4912_/Y _5146_/X _5366_/B vssd1 vssd1 vccd1 vccd1 _5333_/X sky130_fd_sc_hd__o211a_1
X_3594_ _3482_/A _3593_/C _3593_/A vssd1 vssd1 vccd1 vccd1 _3596_/B sky130_fd_sc_hd__a21o_1
X_5264_ _5792_/B vssd1 vssd1 vccd1 vccd1 _5917_/C sky130_fd_sc_hd__clkbuf_4
X_5195_ _5195_/A _5520_/A _5517_/A vssd1 vssd1 vccd1 vccd1 _5196_/B sky130_fd_sc_hd__and3_1
X_4215_ _4516_/C _4209_/B _4219_/A vssd1 vssd1 vccd1 vccd1 _4215_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4146_ _4008_/X _4012_/Y _4138_/Y _4145_/Y vssd1 vssd1 vccd1 vccd1 _4157_/A sky130_fd_sc_hd__o211ai_2
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4077_ _4071_/Y _4073_/Y _3441_/X _5034_/B vssd1 vssd1 vccd1 vccd1 _4284_/A sky130_fd_sc_hd__o2bb2ai_2
XFILLER_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4979_ _4793_/X _4798_/Y _4976_/Y _4978_/Y vssd1 vssd1 vccd1 vccd1 _4979_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4000_ _4160_/A _4160_/B _4160_/C vssd1 vssd1 vccd1 vccd1 _4002_/B sky130_fd_sc_hd__nand3_1
XFILLER_65_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5951_ _5945_/Y _5944_/Y _5943_/Y _5940_/Y vssd1 vssd1 vccd1 vccd1 _5952_/C sky130_fd_sc_hd__o211ai_1
XFILLER_65_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4902_ _4902_/A vssd1 vssd1 vccd1 vccd1 _4903_/B sky130_fd_sc_hd__buf_2
X_5882_ _5872_/Y _5879_/Y _5881_/X vssd1 vssd1 vccd1 vccd1 _5883_/C sky130_fd_sc_hd__a21bo_1
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4833_ _4827_/X _4832_/X _4824_/Y _4819_/Y vssd1 vssd1 vccd1 vccd1 _5190_/B sky130_fd_sc_hd__o211a_1
X_4764_ _4762_/X _4763_/Y _4742_/X _4749_/Y vssd1 vssd1 vccd1 vccd1 _4765_/C sky130_fd_sc_hd__o211ai_1
X_3715_ _4363_/A vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__buf_4
X_4695_ _3448_/X _5446_/A _4529_/B _4932_/A _4694_/X vssd1 vssd1 vccd1 vccd1 _4702_/B
+ sky130_fd_sc_hd__o221ai_4
X_3646_ _5240_/A _4935_/A vssd1 vssd1 vccd1 vccd1 _3646_/Y sky130_fd_sc_hd__nand2_1
X_3577_ _3703_/A _3577_/B _3703_/B vssd1 vssd1 vccd1 vccd1 _3609_/B sky130_fd_sc_hd__nand3_2
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5316_ _5366_/C _5366_/D _5317_/A vssd1 vssd1 vccd1 vccd1 _5316_/Y sky130_fd_sc_hd__a21oi_1
X_6296_ _3310_/A _3190_/C _4832_/C _3190_/A vssd1 vssd1 vccd1 vccd1 _6297_/B sky130_fd_sc_hd__a22oi_2
X_5247_ _5397_/B vssd1 vssd1 vccd1 vccd1 _5918_/B sky130_fd_sc_hd__buf_2
XFILLER_29_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5178_ _5178_/A _5178_/B vssd1 vssd1 vccd1 vccd1 _5178_/Y sky130_fd_sc_hd__nand2_1
X_4129_ _3911_/C _4097_/Y _4128_/Y _4095_/B vssd1 vssd1 vccd1 vccd1 _4130_/B sky130_fd_sc_hd__o211ai_2
XFILLER_56_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3500_ _3500_/A vssd1 vssd1 vccd1 vccd1 _5134_/A sky130_fd_sc_hd__buf_4
X_4480_ _4468_/Y _4469_/Y _4470_/Y _4479_/X vssd1 vssd1 vccd1 vccd1 _4481_/A sky130_fd_sc_hd__o211ai_2
X_3431_ _3766_/A vssd1 vssd1 vccd1 vccd1 _3774_/B sky130_fd_sc_hd__clkbuf_2
X_6150_ _6151_/A _6151_/B _6149_/Y vssd1 vssd1 vccd1 vccd1 _6150_/Y sky130_fd_sc_hd__o21ai_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _4941_/A _5596_/A _5678_/A _3334_/A vssd1 vssd1 vccd1 vccd1 _3362_/Y sky130_fd_sc_hd__a22oi_4
X_5101_ _4922_/A _5100_/A _5100_/B vssd1 vssd1 vccd1 vccd1 _5101_/X sky130_fd_sc_hd__a21o_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6081_ _6081_/A _6081_/B vssd1 vssd1 vccd1 vccd1 _6084_/B sky130_fd_sc_hd__nand2_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3458_/B _4540_/B _4363_/A _3458_/A vssd1 vssd1 vccd1 vccd1 _3293_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_57_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5032_ _5032_/A _5032_/B _5032_/C vssd1 vssd1 vccd1 vccd1 _5310_/A sky130_fd_sc_hd__nand3_2
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5934_ _5933_/A _5933_/B _4287_/B _6171_/C vssd1 vssd1 vccd1 vccd1 _5935_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5865_ _5865_/A _5865_/B _5865_/C vssd1 vssd1 vccd1 vccd1 _5865_/X sky130_fd_sc_hd__and3_1
XFILLER_21_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4816_ _4816_/A vssd1 vssd1 vccd1 vccd1 _4822_/C sky130_fd_sc_hd__buf_2
XFILLER_21_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5796_ _5788_/Y _5790_/X _5791_/Y _5795_/X vssd1 vssd1 vccd1 vccd1 _5823_/A sky130_fd_sc_hd__o211ai_4
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4747_ _4747_/A _6171_/A vssd1 vssd1 vccd1 vccd1 _4748_/B sky130_fd_sc_hd__nor2_1
X_4678_ _4678_/A _4680_/D vssd1 vssd1 vccd1 vccd1 _4679_/A sky130_fd_sc_hd__nand2_1
X_3629_ _4110_/B vssd1 vssd1 vccd1 vccd1 _5834_/A sky130_fd_sc_hd__buf_4
Xoutput49 _5780_/Y vssd1 vssd1 vccd1 vccd1 r[22] sky130_fd_sc_hd__buf_2
Xoutput38 _4168_/Y vssd1 vssd1 vccd1 vccd1 r[12] sky130_fd_sc_hd__buf_2
X_6279_ _6226_/X _6275_/B _6275_/C _6277_/Y _6278_/X vssd1 vssd1 vccd1 vccd1 _6289_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3980_ _3980_/A _3980_/B vssd1 vssd1 vccd1 vccd1 _3980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5650_ _5917_/C vssd1 vssd1 vccd1 vccd1 _6077_/B sky130_fd_sc_hd__clkbuf_2
X_4601_ _4601_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _4601_/Y sky130_fd_sc_hd__nand2_1
X_5581_ _5399_/Y _5580_/Y _5662_/A _5674_/A vssd1 vssd1 vccd1 vccd1 _5585_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4532_ _4532_/A _5539_/A vssd1 vssd1 vccd1 vccd1 _4698_/A sky130_fd_sc_hd__nand2_1
X_4463_ _4463_/A _4463_/B _4463_/C vssd1 vssd1 vccd1 vccd1 _4466_/B sky130_fd_sc_hd__nand3_2
X_6202_ _6202_/A _6202_/B _4830_/A _6244_/A vssd1 vssd1 vccd1 vccd1 _6244_/B sky130_fd_sc_hd__or4bb_2
X_3414_ _3866_/A _3414_/B vssd1 vssd1 vccd1 vccd1 _3552_/A sky130_fd_sc_hd__nand2_2
X_4394_ _4397_/A _4397_/B _4397_/C vssd1 vssd1 vccd1 vccd1 _4394_/X sky130_fd_sc_hd__and3_1
X_6133_ _6132_/Y _6129_/Y _6130_/X vssd1 vssd1 vccd1 vccd1 _6139_/B sky130_fd_sc_hd__a21o_1
X_3345_ _3345_/A _3345_/B vssd1 vssd1 vccd1 vccd1 _3345_/Y sky130_fd_sc_hd__nand2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _3276_/A _3276_/B vssd1 vssd1 vccd1 vccd1 _3287_/A sky130_fd_sc_hd__nand2_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6064_/A _6064_/B vssd1 vssd1 vccd1 vccd1 _6072_/A sky130_fd_sc_hd__nand2_1
X_5015_ _4845_/B _4848_/B _5518_/B vssd1 vssd1 vccd1 vccd1 _5017_/A sky130_fd_sc_hd__a21o_1
XFILLER_38_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5917_ _5917_/A _6009_/A _5917_/C _6002_/B vssd1 vssd1 vccd1 vccd1 _5927_/C sky130_fd_sc_hd__nand4_2
X_5848_ _5914_/B _5843_/Y _5845_/Y _5847_/Y vssd1 vssd1 vccd1 vccd1 _5848_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5779_ _5523_/B _5975_/A _5778_/X vssd1 vssd1 vccd1 vccd1 _5780_/B sky130_fd_sc_hd__o21ai_2
XFILLER_88_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3963_ _4038_/B vssd1 vssd1 vccd1 vccd1 _6010_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5702_ _5542_/B _5793_/A _5809_/A _4179_/X _5799_/A vssd1 vssd1 vccd1 vccd1 _5703_/C
+ sky130_fd_sc_hd__o2111ai_1
X_3894_ _3894_/A _4460_/B vssd1 vssd1 vccd1 vccd1 _3895_/B sky130_fd_sc_hd__nor2_1
X_5633_ _5634_/A _5634_/B _5634_/C _5628_/A vssd1 vssd1 vccd1 vccd1 _5635_/B sky130_fd_sc_hd__a22o_1
X_5564_ _5461_/B _5468_/D _5468_/C vssd1 vssd1 vccd1 vccd1 _5567_/C sky130_fd_sc_hd__a21boi_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4515_ _4681_/A _4681_/B _4508_/Y _4511_/Y vssd1 vssd1 vccd1 vccd1 _4517_/B sky130_fd_sc_hd__o22ai_1
X_5495_ _5495_/A vssd1 vssd1 vccd1 vccd1 _5495_/Y sky130_fd_sc_hd__inv_2
X_4446_ _4436_/Y _4442_/X _4444_/Y _4445_/X vssd1 vssd1 vccd1 vccd1 _4463_/B sky130_fd_sc_hd__o211ai_4
X_4377_ _4564_/A _4564_/B _4564_/C vssd1 vssd1 vccd1 vccd1 _4377_/Y sky130_fd_sc_hd__nand3_2
X_6116_ _5984_/X _6059_/B _6059_/A vssd1 vssd1 vccd1 vccd1 _6116_/X sky130_fd_sc_hd__a21bo_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ input9/X vssd1 vssd1 vccd1 vccd1 _4874_/A sky130_fd_sc_hd__buf_2
XFILLER_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6047_ _6047_/A _6047_/B _6105_/A vssd1 vssd1 vccd1 vccd1 _6048_/B sky130_fd_sc_hd__nand3_1
XFILLER_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3259_ _4540_/A _5251_/A _4235_/B _4355_/B vssd1 vssd1 vccd1 vccd1 _3265_/A sky130_fd_sc_hd__a22o_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5280_ _5281_/A _5281_/B _5219_/X _5220_/Y vssd1 vssd1 vccd1 vccd1 _5427_/A sky130_fd_sc_hd__o2bb2ai_2
X_4300_ _4284_/X _4290_/Y _4298_/Y _4299_/X vssd1 vssd1 vccd1 vccd1 _4308_/B sky130_fd_sc_hd__o211ai_4
XFILLER_4_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4231_ _4239_/A _4239_/B _4230_/Y vssd1 vssd1 vccd1 vccd1 _4231_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4162_ _4166_/B _4165_/A _4160_/X _4161_/Y vssd1 vssd1 vccd1 vccd1 _4338_/A sky130_fd_sc_hd__o2bb2ai_4
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4093_ _4100_/A _4100_/B _4100_/C vssd1 vssd1 vccd1 vccd1 _4095_/B sky130_fd_sc_hd__nand3_4
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4995_ _4995_/A vssd1 vssd1 vccd1 vccd1 _4995_/Y sky130_fd_sc_hd__inv_2
X_3946_ _3946_/A _4133_/A _3984_/C vssd1 vssd1 vccd1 vccd1 _4008_/C sky130_fd_sc_hd__nand3_1
X_3877_ _3787_/B _4103_/A _3803_/B _5401_/A _3868_/Y vssd1 vssd1 vccd1 vccd1 _3878_/B
+ sky130_fd_sc_hd__o2111ai_4
X_5616_ _5616_/A _5616_/B vssd1 vssd1 vccd1 vccd1 _5625_/C sky130_fd_sc_hd__nand2_1
X_5547_ _4080_/X _4363_/D _5704_/A _5794_/A vssd1 vssd1 vccd1 vccd1 _5547_/Y sky130_fd_sc_hd__a22oi_2
X_5478_ _5418_/Y _5426_/Y _5624_/A _5623_/A vssd1 vssd1 vccd1 vccd1 _5483_/B sky130_fd_sc_hd__o211ai_1
X_4429_ _4429_/A _4581_/A vssd1 vssd1 vccd1 vccd1 _4600_/A sky130_fd_sc_hd__nand2_2
XFILLER_86_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3800_ _5209_/A vssd1 vssd1 vccd1 vccd1 _5831_/A sky130_fd_sc_hd__buf_2
X_4780_ _4784_/A _4784_/B _4779_/Y vssd1 vssd1 vccd1 vccd1 _4781_/C sky130_fd_sc_hd__a21o_1
XFILLER_60_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3731_ _3848_/A _3829_/C _3731_/C vssd1 vssd1 vccd1 vccd1 _3845_/B sky130_fd_sc_hd__and3_1
XFILLER_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3662_ _4407_/A vssd1 vssd1 vccd1 vccd1 _4234_/A sky130_fd_sc_hd__clkbuf_2
X_5401_ _5401_/A _5411_/C vssd1 vssd1 vccd1 vccd1 _5402_/B sky130_fd_sc_hd__nand2_1
X_3593_ _3593_/A _3593_/B _3593_/C vssd1 vssd1 vccd1 vccd1 _3596_/A sky130_fd_sc_hd__nand3_1
X_5332_ _5337_/A _5332_/B vssd1 vssd1 vccd1 vccd1 _5335_/A sky130_fd_sc_hd__nand2_1
X_5263_ _5263_/A _5263_/B _5263_/C _6010_/B vssd1 vssd1 vccd1 vccd1 _5420_/B sky130_fd_sc_hd__nand4_4
X_5194_ _5517_/A _5520_/A _5195_/A vssd1 vssd1 vccd1 vccd1 _5196_/A sky130_fd_sc_hd__a21oi_1
X_4214_ _4194_/Y _4198_/Y _4213_/Y vssd1 vssd1 vccd1 vccd1 _4219_/A sky130_fd_sc_hd__o21ai_1
X_4145_ _4317_/A _4141_/Y _4142_/Y _4144_/X vssd1 vssd1 vccd1 vccd1 _4145_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4076_ _4777_/D vssd1 vssd1 vccd1 vccd1 _5034_/B sky130_fd_sc_hd__inv_4
XFILLER_83_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4978_ _4643_/B _4795_/Y _4977_/Y _4797_/Y vssd1 vssd1 vccd1 vccd1 _4978_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3929_ _3945_/A vssd1 vssd1 vccd1 vccd1 _3929_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5950_ _5816_/B _5822_/Y _5940_/Y _5943_/Y vssd1 vssd1 vccd1 vccd1 _5952_/B sky130_fd_sc_hd__a22o_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4901_ _4901_/A _4901_/B vssd1 vssd1 vccd1 vccd1 _4902_/A sky130_fd_sc_hd__nand2_1
X_5881_ _5556_/Y _5694_/X _5750_/Y _5723_/Y vssd1 vssd1 vccd1 vccd1 _5881_/X sky130_fd_sc_hd__o31a_1
X_4832_ _4832_/A _6255_/B _4832_/C vssd1 vssd1 vccd1 vccd1 _4832_/X sky130_fd_sc_hd__and3_1
XFILLER_60_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4763_ _4890_/A _4890_/B _4762_/A vssd1 vssd1 vccd1 vccd1 _4763_/Y sky130_fd_sc_hd__a21oi_1
X_3714_ _5596_/A _5596_/B _5132_/A _3714_/D vssd1 vssd1 vccd1 vccd1 _3714_/X sky130_fd_sc_hd__and4_1
X_4694_ _5299_/B _5696_/A _5284_/D _3543_/B vssd1 vssd1 vccd1 vccd1 _4694_/X sky130_fd_sc_hd__a22o_1
X_3645_ _3758_/B vssd1 vssd1 vccd1 vccd1 _4935_/A sky130_fd_sc_hd__buf_2
X_3576_ _3576_/A _3730_/B vssd1 vssd1 vccd1 vccd1 _3703_/A sky130_fd_sc_hd__nand2_1
X_5315_ _5130_/C _5130_/A _5130_/B _5142_/X vssd1 vssd1 vccd1 vccd1 _5317_/A sky130_fd_sc_hd__a31oi_2
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6295_ _6295_/A _6295_/B vssd1 vssd1 vccd1 vccd1 _6295_/X sky130_fd_sc_hd__xor2_4
X_5246_ _5250_/B vssd1 vssd1 vccd1 vccd1 _5246_/X sky130_fd_sc_hd__buf_4
X_5177_ _5177_/A vssd1 vssd1 vccd1 vccd1 _5177_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4128_ _4128_/A _4128_/B vssd1 vssd1 vccd1 vccd1 _4128_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4059_ _4868_/A _4777_/D vssd1 vssd1 vccd1 vccd1 _4059_/Y sky130_fd_sc_hd__nand2_2
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3430_ _4730_/A vssd1 vssd1 vccd1 vccd1 _4571_/A sky130_fd_sc_hd__buf_2
X_3361_ _3344_/Y _3349_/Y _3477_/A vssd1 vssd1 vccd1 vccd1 _3372_/A sky130_fd_sc_hd__o21ai_1
X_6080_ _6081_/A _6081_/B _6084_/A vssd1 vssd1 vccd1 vccd1 _6087_/A sky130_fd_sc_hd__a21o_1
X_5100_ _5100_/A _5100_/B vssd1 vssd1 vccd1 vccd1 _5100_/Y sky130_fd_sc_hd__nand2_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _4903_/B _5208_/A _5582_/A _5805_/A _5025_/Y vssd1 vssd1 vccd1 vccd1 _5032_/C
+ sky130_fd_sc_hd__o2111ai_4
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _3533_/A vssd1 vssd1 vccd1 vccd1 _3458_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5933_ _5933_/A _5933_/B _5933_/C _5933_/D vssd1 vssd1 vccd1 vccd1 _5935_/A sky130_fd_sc_hd__and4_1
X_5864_ _5957_/B _5829_/X _5859_/Y _5860_/Y _5863_/X vssd1 vssd1 vccd1 vccd1 _5872_/B
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_61_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4815_ _4815_/A _4815_/B _4815_/C vssd1 vssd1 vccd1 vccd1 _4816_/A sky130_fd_sc_hd__nand3_1
X_5795_ _4179_/X _5407_/C _5793_/Y _5794_/Y vssd1 vssd1 vccd1 vccd1 _5795_/X sky130_fd_sc_hd__a22o_1
X_4746_ _4746_/A _4746_/B vssd1 vssd1 vccd1 vccd1 _4748_/A sky130_fd_sc_hd__nand2_1
X_4677_ _4508_/Y _4525_/X _4672_/Y _4676_/X vssd1 vssd1 vccd1 vccd1 _4842_/C sky130_fd_sc_hd__o211ai_2
X_3628_ _5212_/A vssd1 vssd1 vccd1 vccd1 _4110_/B sky130_fd_sc_hd__buf_2
Xoutput39 _4342_/X vssd1 vssd1 vccd1 vccd1 r[13] sky130_fd_sc_hd__buf_2
X_3559_ _3559_/A _3559_/B vssd1 vssd1 vccd1 vccd1 _3560_/B sky130_fd_sc_hd__nand2_2
X_6278_ _6266_/A _6266_/B _6266_/C _6247_/B _6247_/A vssd1 vssd1 vccd1 vccd1 _6278_/X
+ sky130_fd_sc_hd__a311o_1
X_5229_ _5229_/A _5240_/D vssd1 vssd1 vccd1 vccd1 _5229_/Y sky130_fd_sc_hd__nand2_2
XFILLER_29_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4600_ _4600_/A _4600_/B _4600_/C vssd1 vssd1 vccd1 vccd1 _4600_/X sky130_fd_sc_hd__and3_1
XFILLER_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5580_ _5580_/A _5919_/B vssd1 vssd1 vccd1 vccd1 _5580_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4531_ _4363_/A _5553_/B _4529_/Y _4530_/Y vssd1 vssd1 vccd1 vccd1 _4531_/Y sky130_fd_sc_hd__a22oi_4
X_4462_ _4453_/Y _4459_/Y _4461_/Y vssd1 vssd1 vccd1 vccd1 _4463_/C sky130_fd_sc_hd__o21ai_2
X_6201_ _6233_/A _6233_/B _6203_/C _6233_/C vssd1 vssd1 vccd1 vccd1 _6244_/A sky130_fd_sc_hd__nand4_2
X_3413_ _4460_/A vssd1 vssd1 vccd1 vccd1 _3474_/A sky130_fd_sc_hd__buf_4
X_4393_ _4367_/Y _4371_/Y _4377_/Y _4392_/Y vssd1 vssd1 vccd1 vccd1 _4397_/C sky130_fd_sc_hd__o211ai_4
X_6132_ _6132_/A _6132_/B _6132_/C _6170_/D vssd1 vssd1 vccd1 vccd1 _6132_/Y sky130_fd_sc_hd__nand4_2
X_3344_ _3358_/D _3440_/A _3348_/A vssd1 vssd1 vccd1 vccd1 _3344_/Y sky130_fd_sc_hd__a21oi_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3275_ _4432_/A _3870_/A vssd1 vssd1 vccd1 vccd1 _3276_/B sky130_fd_sc_hd__nand2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6127_/A _6127_/C vssd1 vssd1 vccd1 vccd1 _6064_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5014_ _5014_/A _5014_/B vssd1 vssd1 vccd1 vccd1 _5518_/B sky130_fd_sc_hd__nand2_2
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5916_ _6010_/A vssd1 vssd1 vccd1 vccd1 _6132_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_41_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5847_ _5847_/A _5847_/B vssd1 vssd1 vccd1 vccd1 _5847_/Y sky130_fd_sc_hd__nand2_1
X_5778_ _5776_/A _5776_/C _5777_/Y vssd1 vssd1 vccd1 vccd1 _5778_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4729_ _4729_/A vssd1 vssd1 vccd1 vccd1 _4809_/B sky130_fd_sc_hd__buf_2
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5701_ _5701_/A _5701_/B vssd1 vssd1 vccd1 vccd1 _5793_/A sky130_fd_sc_hd__nand2_1
X_3962_ _4936_/B vssd1 vssd1 vccd1 vccd1 _4038_/B sky130_fd_sc_hd__buf_2
X_3893_ _3891_/A _4064_/A _3889_/A _3747_/B vssd1 vssd1 vccd1 vccd1 _3895_/A sky130_fd_sc_hd__o2bb2ai_1
X_5632_ _5502_/A _5502_/C _5525_/A vssd1 vssd1 vccd1 vccd1 _5635_/A sky130_fd_sc_hd__a21boi_2
X_5563_ _5563_/A _5563_/B _5563_/C vssd1 vssd1 vccd1 vccd1 _5567_/B sky130_fd_sc_hd__nand3_1
X_4514_ _4519_/B _4514_/B _4514_/C vssd1 vssd1 vccd1 vccd1 _4842_/A sky130_fd_sc_hd__nand3_1
X_5494_ _5494_/A vssd1 vssd1 vccd1 vccd1 _5525_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4445_ _4600_/A _4600_/B _4443_/Y vssd1 vssd1 vccd1 vccd1 _4445_/X sky130_fd_sc_hd__a21o_1
X_4376_ _4197_/A _4196_/Y _4197_/B vssd1 vssd1 vccd1 vccd1 _4564_/C sky130_fd_sc_hd__o21ai_4
X_6115_ _6193_/A _6193_/B vssd1 vssd1 vccd1 vccd1 _6220_/A sky130_fd_sc_hd__nor2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _4355_/B vssd1 vssd1 vccd1 vccd1 _4542_/A sky130_fd_sc_hd__clkbuf_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6046_ _6047_/A _6047_/B _6105_/A vssd1 vssd1 vccd1 vccd1 _6048_/A sky130_fd_sc_hd__a21o_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _4877_/A vssd1 vssd1 vccd1 vccd1 _5251_/A sky130_fd_sc_hd__clkbuf_4
X_3189_ _3189_/A vssd1 vssd1 vccd1 vccd1 _5603_/A sky130_fd_sc_hd__buf_4
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4230_ _4530_/A _5037_/A vssd1 vssd1 vccd1 vccd1 _4230_/Y sky130_fd_sc_hd__nand2_2
X_4161_ _4161_/A _4161_/B vssd1 vssd1 vccd1 vccd1 _4161_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4092_ _4100_/A _4100_/B _4100_/C vssd1 vssd1 vccd1 vccd1 _4095_/A sky130_fd_sc_hd__a21o_1
XFILLER_67_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4994_ _4986_/X _4991_/Y _5021_/A vssd1 vssd1 vccd1 vccd1 _5020_/A sky130_fd_sc_hd__o21bai_1
X_3945_ _3945_/A vssd1 vssd1 vccd1 vccd1 _4133_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5615_ _5612_/X _5613_/Y _5614_/Y vssd1 vssd1 vccd1 vccd1 _5616_/B sky130_fd_sc_hd__o21ai_1
X_3876_ _3868_/Y _3872_/Y _3873_/Y vssd1 vssd1 vccd1 vccd1 _3878_/A sky130_fd_sc_hd__a21bo_1
X_5546_ _5546_/A _5925_/A vssd1 vssd1 vccd1 vccd1 _5546_/Y sky130_fd_sc_hd__nand2_1
X_5477_ _5477_/A _5477_/B vssd1 vssd1 vccd1 vccd1 _5623_/A sky130_fd_sc_hd__nand2_1
X_4428_ _5045_/A _4877_/D vssd1 vssd1 vccd1 vccd1 _4581_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4359_ _4680_/A _4362_/B _3186_/X _6171_/C vssd1 vssd1 vccd1 vccd1 _4359_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_86_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ _6091_/A _6091_/B _6027_/X vssd1 vssd1 vccd1 vccd1 _6030_/B sky130_fd_sc_hd__a21o_1
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3730_ _3730_/A _3730_/B vssd1 vssd1 vccd1 vccd1 _3848_/A sky130_fd_sc_hd__nand2_1
X_3661_ _3903_/A vssd1 vssd1 vccd1 vccd1 _4930_/A sky130_fd_sc_hd__buf_2
X_5400_ _5403_/A _5674_/A _5399_/Y _5208_/B vssd1 vssd1 vccd1 vccd1 _5402_/A sky130_fd_sc_hd__o2bb2ai_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3592_ _3592_/A vssd1 vssd1 vccd1 vccd1 _3593_/A sky130_fd_sc_hd__inv_2
X_5331_ _5331_/A _5331_/B _5331_/C vssd1 vssd1 vccd1 vccd1 _5332_/B sky130_fd_sc_hd__nand3_1
X_5262_ _5792_/B vssd1 vssd1 vccd1 vccd1 _6010_/B sky130_fd_sc_hd__clkbuf_4
X_5193_ _5518_/A _5518_/B _4847_/B _5192_/Y vssd1 vssd1 vccd1 vccd1 _5195_/A sky130_fd_sc_hd__o31a_1
XFILLER_68_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4213_ _4213_/A _4213_/B _4213_/C vssd1 vssd1 vccd1 vccd1 _4213_/Y sky130_fd_sc_hd__nand3_2
X_4144_ _3968_/A _4143_/X _4044_/A _4051_/A vssd1 vssd1 vccd1 vccd1 _4144_/X sky130_fd_sc_hd__o211a_1
X_4075_ _4060_/Y _4063_/Y _4070_/X _4074_/X vssd1 vssd1 vccd1 vccd1 _4100_/A sky130_fd_sc_hd__o211ai_4
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4977_ _4801_/A _4801_/B _4796_/A _4796_/B vssd1 vssd1 vccd1 vccd1 _4977_/Y sky130_fd_sc_hd__o2bb2ai_1
X_3928_ _3928_/A _3928_/B _3928_/C vssd1 vssd1 vccd1 vccd1 _3945_/A sky130_fd_sc_hd__nand3_2
X_3859_ _3859_/A _3859_/B vssd1 vssd1 vccd1 vccd1 _3859_/X sky130_fd_sc_hd__xor2_2
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5529_ _5623_/A _5528_/Y _5623_/B vssd1 vssd1 vccd1 vccd1 _5622_/A sky130_fd_sc_hd__o21ai_1
XFILLER_59_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5880_ _5748_/X _5740_/X _5872_/Y _5879_/Y vssd1 vssd1 vccd1 vccd1 _5883_/B sky130_fd_sc_hd__o211ai_2
XFILLER_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4900_ _4904_/B _5284_/C vssd1 vssd1 vccd1 vccd1 _4903_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4831_ _5352_/A vssd1 vssd1 vccd1 vccd1 _6255_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4762_ _4762_/A _4890_/A _4890_/B vssd1 vssd1 vccd1 vccd1 _4762_/X sky130_fd_sc_hd__and3_1
X_3713_ _5372_/B _4363_/B _3714_/D _3677_/A vssd1 vssd1 vccd1 vccd1 _3713_/Y sky130_fd_sc_hd__a22oi_2
X_4693_ _4693_/A _5119_/D vssd1 vssd1 vccd1 vccd1 _4932_/A sky130_fd_sc_hd__nand2_4
X_3644_ _3558_/A _3560_/B _3565_/Y _3564_/X vssd1 vssd1 vccd1 vccd1 _3689_/A sky130_fd_sc_hd__o2bb2ai_2
XFILLER_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3575_ _3570_/Y _3478_/A _3486_/C vssd1 vssd1 vccd1 vccd1 _3575_/Y sky130_fd_sc_hd__a21oi_1
X_5314_ _5321_/C vssd1 vssd1 vccd1 vccd1 _5366_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6294_ _6294_/A _6294_/B _6294_/C vssd1 vssd1 vccd1 vccd1 _6295_/B sky130_fd_sc_hd__and3_1
X_5245_ _5245_/A _5245_/B vssd1 vssd1 vccd1 vccd1 _5250_/B sky130_fd_sc_hd__nand2_2
X_5176_ _5176_/A _5176_/B vssd1 vssd1 vccd1 vccd1 _5180_/B sky130_fd_sc_hd__nand2_1
X_4127_ _4135_/C _4135_/B _4127_/C vssd1 vssd1 vccd1 vccd1 _4127_/X sky130_fd_sc_hd__and3_1
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4058_ _4065_/A vssd1 vssd1 vccd1 vccd1 _4777_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3360_ _3360_/A vssd1 vssd1 vccd1 vccd1 _3477_/A sky130_fd_sc_hd__clkbuf_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5284_/C vssd1 vssd1 vccd1 vccd1 _5805_/A sky130_fd_sc_hd__clkbuf_4
X_3291_ _4730_/A vssd1 vssd1 vccd1 vccd1 _3533_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_78_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5932_ _6020_/C _6079_/A _6077_/A _6076_/B vssd1 vssd1 vccd1 vccd1 _5933_/B sky130_fd_sc_hd__nand4_4
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5863_ _5957_/A _5865_/B _5865_/C vssd1 vssd1 vccd1 vccd1 _5863_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5794_ _5794_/A _5794_/B _5794_/C _5918_/B vssd1 vssd1 vccd1 vccd1 _5794_/Y sky130_fd_sc_hd__nand4_1
X_4814_ _4814_/A _4814_/B vssd1 vssd1 vccd1 vccd1 _4815_/C sky130_fd_sc_hd__nand2_1
XFILLER_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4745_ _4745_/A _4746_/A _4746_/B vssd1 vssd1 vccd1 vccd1 _4745_/Y sky130_fd_sc_hd__nand3_2
X_4676_ _4680_/C _4680_/D _4679_/B vssd1 vssd1 vccd1 vccd1 _4676_/X sky130_fd_sc_hd__a21o_1
X_3627_ _3617_/A _3630_/B _3626_/X vssd1 vssd1 vccd1 vccd1 _3632_/A sky130_fd_sc_hd__a21o_1
X_3558_ _3558_/A _3558_/B vssd1 vssd1 vccd1 vccd1 _3560_/A sky130_fd_sc_hd__nand2_1
X_6277_ _6277_/A vssd1 vssd1 vccd1 vccd1 _6277_/Y sky130_fd_sc_hd__inv_2
X_3489_ _3510_/A vssd1 vssd1 vccd1 vccd1 _5212_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5228_ _5095_/B _5227_/Y _5095_/A vssd1 vssd1 vccd1 vccd1 _5256_/A sky130_fd_sc_hd__a21boi_4
X_5159_ _5159_/A _5159_/B _5159_/C vssd1 vssd1 vccd1 vccd1 _5171_/C sky130_fd_sc_hd__nand3_2
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4530_ _4530_/A _4945_/A _4530_/C _5284_/D vssd1 vssd1 vccd1 vccd1 _4530_/Y sky130_fd_sc_hd__nand4_2
XFILLER_7_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4461_ _4476_/A _4461_/B vssd1 vssd1 vccd1 vccd1 _4461_/Y sky130_fd_sc_hd__nand2_1
X_6200_ _6233_/B _6203_/C _6233_/C _6233_/A vssd1 vssd1 vccd1 vccd1 _6202_/A sky130_fd_sc_hd__a22oi_1
X_3412_ _4025_/A vssd1 vssd1 vccd1 vccd1 _3468_/A sky130_fd_sc_hd__clkinv_2
X_6131_ _6235_/B _6128_/Y _6129_/Y _6130_/X vssd1 vssd1 vccd1 vccd1 _6131_/X sky130_fd_sc_hd__o211a_1
X_4392_ _4386_/Y _4680_/B _4391_/X vssd1 vssd1 vccd1 vccd1 _4392_/Y sky130_fd_sc_hd__o21ai_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _5231_/A _3500_/A vssd1 vssd1 vccd1 vccd1 _3348_/A sky130_fd_sc_hd__nand2_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _4730_/A vssd1 vssd1 vccd1 vccd1 _4432_/A sky130_fd_sc_hd__buf_4
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6127_/B _6065_/C vssd1 vssd1 vccd1 vccd1 _6064_/A sky130_fd_sc_hd__nand2_1
X_5013_ _5012_/B _5012_/C _5012_/A vssd1 vssd1 vccd1 vccd1 _5014_/B sky130_fd_sc_hd__a21o_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5915_ _5868_/A _5868_/B _5868_/C _5989_/A _6024_/A vssd1 vssd1 vccd1 vccd1 _5949_/B
+ sky130_fd_sc_hd__a32o_1
X_5846_ _5846_/A _5846_/B vssd1 vssd1 vccd1 vccd1 _5847_/A sky130_fd_sc_hd__nand2_1
X_5777_ _5639_/B _5639_/C _5639_/A vssd1 vssd1 vccd1 vccd1 _5777_/Y sky130_fd_sc_hd__a21oi_1
X_4728_ _4975_/A _4975_/B _4975_/C vssd1 vssd1 vccd1 vccd1 _4729_/A sky130_fd_sc_hd__and3_1
X_4659_ _4659_/A _4659_/B vssd1 vssd1 vccd1 vccd1 _4660_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3961_ _3521_/A _6165_/B _3964_/A _3964_/B vssd1 vssd1 vccd1 vccd1 _4143_/A sky130_fd_sc_hd__a22oi_4
X_5700_ _5554_/B _5542_/Y _5540_/X _5538_/X vssd1 vssd1 vccd1 vccd1 _5703_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_16_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3892_ _3894_/A _4460_/B _3747_/B _4071_/A _3891_/Y vssd1 vssd1 vccd1 vccd1 _4097_/A
+ sky130_fd_sc_hd__o221ai_4
X_5631_ _5631_/A _5631_/B _5631_/C vssd1 vssd1 vccd1 vccd1 _5640_/C sky130_fd_sc_hd__nand3_2
X_5562_ _5413_/B _5413_/C _5414_/Y vssd1 vssd1 vccd1 vccd1 _5563_/C sky130_fd_sc_hd__a21o_1
X_4513_ _4519_/B _4514_/B _4514_/C vssd1 vssd1 vccd1 vccd1 _4513_/X sky130_fd_sc_hd__and3_1
X_5493_ _5493_/A _5493_/B _5493_/C vssd1 vssd1 vccd1 vccd1 _5494_/A sky130_fd_sc_hd__nand3_1
XFILLER_7_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4444_ _4267_/Y _4568_/A _4600_/A _4443_/Y vssd1 vssd1 vccd1 vccd1 _4444_/Y sky130_fd_sc_hd__o211ai_2
X_4375_ _4182_/B _4529_/A _4941_/A _4186_/B _4365_/Y vssd1 vssd1 vccd1 vccd1 _4564_/B
+ sky130_fd_sc_hd__o2111ai_4
X_6114_ _6219_/C _6219_/B vssd1 vssd1 vccd1 vccd1 _6118_/A sky130_fd_sc_hd__nand2_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _4714_/A vssd1 vssd1 vccd1 vccd1 _3334_/A sky130_fd_sc_hd__buf_4
XFILLER_85_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6045_ _6043_/Y _5943_/B _5940_/Y _6044_/Y vssd1 vssd1 vccd1 vccd1 _6105_/A sky130_fd_sc_hd__a22o_1
XFILLER_58_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3772_/A vssd1 vssd1 vccd1 vccd1 _4877_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3188_ _3441_/A vssd1 vssd1 vccd1 vccd1 _3189_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5829_ _5822_/Y _5944_/B _5827_/Y _5828_/X vssd1 vssd1 vccd1 vccd1 _5829_/X sky130_fd_sc_hd__o211a_1
XFILLER_22_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4160_ _4160_/A _4160_/B _4160_/C vssd1 vssd1 vccd1 vccd1 _4160_/X sky130_fd_sc_hd__and3_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4091_ _4091_/A _4091_/B vssd1 vssd1 vccd1 vccd1 _4100_/C sky130_fd_sc_hd__nand2_2
XFILLER_95_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4993_ _5004_/B vssd1 vssd1 vccd1 vccd1 _5021_/A sky130_fd_sc_hd__inv_2
X_3944_ _3822_/C _3934_/Y _3942_/X _3943_/X vssd1 vssd1 vccd1 vccd1 _4008_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_23_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3875_ _3878_/C _3875_/B _3875_/C vssd1 vssd1 vccd1 vccd1 _3980_/B sky130_fd_sc_hd__nand3b_2
X_5614_ _5614_/A _5614_/B _5614_/C vssd1 vssd1 vccd1 vccd1 _5614_/Y sky130_fd_sc_hd__nand3_4
X_5545_ _5538_/X _5540_/X _5808_/A _4179_/X _5542_/Y vssd1 vssd1 vccd1 vccd1 _5549_/B
+ sky130_fd_sc_hd__o2111ai_4
X_5476_ _5479_/A _5634_/A _5479_/B vssd1 vssd1 vccd1 vccd1 _5477_/B sky130_fd_sc_hd__nand3_1
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4427_ _4569_/A vssd1 vssd1 vccd1 vccd1 _4877_/D sky130_fd_sc_hd__buf_2
XFILLER_48_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ _4387_/A vssd1 vssd1 vccd1 vccd1 _6171_/C sky130_fd_sc_hd__buf_4
X_4289_ _4071_/A _4057_/X _4060_/Y vssd1 vssd1 vccd1 vccd1 _4289_/X sky130_fd_sc_hd__a21o_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _3309_/A _3309_/B _3309_/C vssd1 vssd1 vccd1 vccd1 _3392_/A sky130_fd_sc_hd__nand3_2
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6028_ _6091_/A _6091_/B _6027_/X _6024_/A vssd1 vssd1 vccd1 vccd1 _6030_/A sky130_fd_sc_hd__a31oi_1
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3660_ input7/X vssd1 vssd1 vccd1 vccd1 _4855_/B sky130_fd_sc_hd__buf_2
X_3591_ _3591_/A _3591_/B _3857_/C vssd1 vssd1 vccd1 vccd1 _6294_/A sky130_fd_sc_hd__nand3_2
X_5330_ _5327_/Y _5495_/A _5329_/X _5277_/Y _5283_/Y vssd1 vssd1 vccd1 vccd1 _5331_/C
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5261_ _5082_/Y _5081_/X _5257_/Y _5260_/Y vssd1 vssd1 vccd1 vccd1 _5269_/A sky130_fd_sc_hd__o22ai_4
X_4212_ _4220_/A _4220_/B vssd1 vssd1 vccd1 vccd1 _4212_/Y sky130_fd_sc_hd__nand2_1
X_5192_ _5190_/Y _5014_/A _4839_/A _5191_/Y vssd1 vssd1 vccd1 vccd1 _5192_/Y sky130_fd_sc_hd__a31oi_4
X_4143_ _4143_/A _4143_/B vssd1 vssd1 vccd1 vccd1 _4143_/X sky130_fd_sc_hd__or2_1
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4074_ _4071_/Y _4073_/Y _4059_/Y vssd1 vssd1 vccd1 vccd1 _4074_/X sky130_fd_sc_hd__a21o_1
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4976_ _4976_/A _4976_/B vssd1 vssd1 vccd1 vccd1 _4976_/Y sky130_fd_sc_hd__nand2_2
X_3927_ _3927_/A _4128_/B _3927_/C vssd1 vssd1 vccd1 vccd1 _3928_/C sky130_fd_sc_hd__nand3_1
X_3858_ _3856_/Y _3857_/X _3745_/B _3745_/A vssd1 vssd1 vccd1 vccd1 _3859_/B sky130_fd_sc_hd__a22oi_4
X_3789_ _4026_/A _3866_/A _5655_/A _4904_/B vssd1 vssd1 vccd1 vccd1 _3790_/A sky130_fd_sc_hd__nand4_1
X_5528_ _5490_/A _5490_/B _5490_/C _5490_/D vssd1 vssd1 vccd1 vccd1 _5528_/Y sky130_fd_sc_hd__a22oi_1
X_5459_ _5468_/C _5468_/D vssd1 vssd1 vccd1 vccd1 _5461_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4830_ _4830_/A vssd1 vssd1 vccd1 vccd1 _5352_/A sky130_fd_sc_hd__buf_2
XFILLER_33_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4761_ _4880_/A _4761_/B vssd1 vssd1 vccd1 vccd1 _4762_/A sky130_fd_sc_hd__nand2_1
X_3712_ _4936_/A vssd1 vssd1 vccd1 vccd1 _3714_/D sky130_fd_sc_hd__clkbuf_4
X_4692_ _4365_/B _4533_/X _4690_/Y _4691_/Y vssd1 vssd1 vccd1 vccd1 _4702_/A sky130_fd_sc_hd__o22a_1
X_3643_ _3720_/A _3720_/B vssd1 vssd1 vccd1 vccd1 _3687_/A sky130_fd_sc_hd__nand2_2
X_5313_ _5313_/A _5313_/B _5313_/C vssd1 vssd1 vccd1 vccd1 _5321_/C sky130_fd_sc_hd__nand3_1
X_3574_ _3574_/A _3574_/B _3574_/C vssd1 vssd1 vccd1 vccd1 _3574_/X sky130_fd_sc_hd__and3_1
X_6293_ _3591_/A _3591_/B _3597_/Y vssd1 vssd1 vccd1 vccd1 _6294_/C sky130_fd_sc_hd__a21o_1
X_5244_ _5372_/B _5575_/B _5372_/C _3677_/A vssd1 vssd1 vccd1 vccd1 _5244_/Y sky130_fd_sc_hd__a22oi_4
X_5175_ _5175_/A _5175_/B vssd1 vssd1 vccd1 vccd1 _5176_/B sky130_fd_sc_hd__and2_1
XFILLER_29_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4126_ _4220_/A _4135_/B _4127_/C vssd1 vssd1 vccd1 vccd1 _4126_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4057_ _4071_/B vssd1 vssd1 vccd1 vccd1 _4057_/X sky130_fd_sc_hd__buf_2
XFILLER_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4959_ _4958_/X _4955_/Y _4956_/X vssd1 vssd1 vccd1 vccd1 _4959_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _3500_/A vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__buf_4
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5931_ _5931_/A vssd1 vssd1 vccd1 vccd1 _6079_/A sky130_fd_sc_hd__buf_2
XFILLER_18_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5862_ _5865_/A vssd1 vssd1 vccd1 vccd1 _5957_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5793_ _5793_/A _5793_/B vssd1 vssd1 vccd1 vccd1 _5793_/Y sky130_fd_sc_hd__nand2_1
X_4813_ _4793_/X _4798_/Y _4809_/A _4809_/B _4803_/Y vssd1 vssd1 vccd1 vccd1 _4815_/B
+ sky130_fd_sc_hd__o221ai_1
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4744_ _4744_/A _4877_/D vssd1 vssd1 vccd1 vccd1 _4745_/A sky130_fd_sc_hd__nand2_2
X_4675_ _3186_/X _4674_/X _4386_/Y _4362_/B vssd1 vssd1 vccd1 vccd1 _4679_/B sky130_fd_sc_hd__o31a_2
X_3626_ _4355_/B _4779_/B vssd1 vssd1 vccd1 vccd1 _3626_/X sky130_fd_sc_hd__and2_1
X_3557_ _3558_/A _3558_/B _3559_/A _3559_/B vssd1 vssd1 vccd1 vccd1 _3702_/A sky130_fd_sc_hd__nand4_2
X_6276_ _6195_/Y _6221_/Y _6274_/Y _6275_/Y vssd1 vssd1 vccd1 vccd1 _6289_/B sky130_fd_sc_hd__o211ai_1
X_5227_ _5070_/C _5093_/Y _5078_/Y vssd1 vssd1 vccd1 vccd1 _5227_/Y sky130_fd_sc_hd__a21oi_1
X_3488_ _3584_/C _3584_/A _3584_/B _3592_/A vssd1 vssd1 vccd1 vccd1 _3488_/X sky130_fd_sc_hd__a31o_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5158_ _4989_/Y _4972_/Y _4927_/Y vssd1 vssd1 vccd1 vccd1 _5159_/C sky130_fd_sc_hd__a21oi_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4109_ _3714_/D _5831_/A _5669_/A _5302_/C vssd1 vssd1 vccd1 vccd1 _4109_/Y sky130_fd_sc_hd__a22oi_4
X_5089_ _4871_/A _5075_/Y _5087_/X _5088_/Y vssd1 vssd1 vccd1 vccd1 _5096_/A sky130_fd_sc_hd__o2bb2ai_1
XFILLER_56_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4460_ _4460_/A _4460_/B vssd1 vssd1 vccd1 vccd1 _4461_/B sky130_fd_sc_hd__nor2_1
X_4391_ _4680_/A _4356_/A _4390_/Y vssd1 vssd1 vccd1 vccd1 _4391_/X sky130_fd_sc_hd__a21o_1
X_3411_ _3486_/C vssd1 vssd1 vccd1 vccd1 _3479_/A sky130_fd_sc_hd__inv_2
X_3342_ _3342_/A _3342_/B vssd1 vssd1 vccd1 vccd1 _3440_/A sky130_fd_sc_hd__nand2_2
X_6130_ _6072_/A _6068_/B _6072_/B vssd1 vssd1 vccd1 vccd1 _6130_/X sky130_fd_sc_hd__a21bo_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _5998_/A _5998_/B _5996_/B vssd1 vssd1 vccd1 vccd1 _6061_/X sky130_fd_sc_hd__a21o_1
XFILLER_58_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3273_ input1/X vssd1 vssd1 vccd1 vccd1 _4730_/A sky130_fd_sc_hd__clkbuf_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5012_/A _5012_/B _5012_/C vssd1 vssd1 vccd1 vccd1 _5014_/A sky130_fd_sc_hd__nand3_2
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5914_ _5914_/A _5914_/B _5914_/C _5914_/D vssd1 vssd1 vccd1 vccd1 _6024_/A sky130_fd_sc_hd__nand4_2
X_5845_ _5845_/A _5858_/C _6203_/D _6165_/D vssd1 vssd1 vccd1 vccd1 _5845_/Y sky130_fd_sc_hd__nand4_1
X_5776_ _5776_/A _5776_/B _5776_/C _5776_/D vssd1 vssd1 vccd1 vccd1 _5975_/A sky130_fd_sc_hd__nand4_2
X_4727_ _4689_/B _4689_/A _4549_/X vssd1 vssd1 vccd1 vccd1 _4975_/C sky130_fd_sc_hd__a21oi_1
X_4658_ _4649_/Y _4650_/Y _4645_/Y vssd1 vssd1 vccd1 vccd1 _4660_/A sky130_fd_sc_hd__o21ai_1
X_3609_ _3609_/A _3609_/B _3609_/C vssd1 vssd1 vccd1 vccd1 _3609_/X sky130_fd_sc_hd__and3_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4589_ _5378_/A _5212_/B _5541_/B _3551_/A vssd1 vssd1 vccd1 vccd1 _4589_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6259_ _6260_/A _6260_/B _6258_/A vssd1 vssd1 vccd1 vccd1 _6259_/X sky130_fd_sc_hd__or3b_1
XFILLER_67_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3960_ _4355_/A _3960_/B _5792_/A _4363_/D vssd1 vssd1 vccd1 vccd1 _3964_/B sky130_fd_sc_hd__nand4_4
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3891_ _3891_/A _4064_/A vssd1 vssd1 vccd1 vccd1 _3891_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5630_ _5634_/C _5634_/D _5629_/A vssd1 vssd1 vccd1 vccd1 _5631_/C sky130_fd_sc_hd__a21o_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5561_ _5694_/A _5694_/B _5561_/C _5694_/C vssd1 vssd1 vccd1 vccd1 _5563_/B sky130_fd_sc_hd__nand4_1
X_5492_ _5623_/A _5492_/B vssd1 vssd1 vccd1 vccd1 _5493_/C sky130_fd_sc_hd__nand2_1
X_4512_ _4508_/Y _4511_/Y _4516_/C vssd1 vssd1 vccd1 vccd1 _4514_/C sky130_fd_sc_hd__o21ai_1
X_4443_ _4868_/A _4884_/B vssd1 vssd1 vccd1 vccd1 _4443_/Y sky130_fd_sc_hd__nand2_2
X_4374_ _4363_/Y _4365_/Y _3280_/X _5453_/B vssd1 vssd1 vccd1 vccd1 _4564_/A sky130_fd_sc_hd__o2bb2ai_2
X_6113_ _6112_/A _6112_/B _6112_/C vssd1 vssd1 vccd1 vccd1 _6219_/B sky130_fd_sc_hd__a21o_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _5248_/A vssd1 vssd1 vccd1 vccd1 _5678_/B sky130_fd_sc_hd__buf_4
X_6044_ _5816_/A _5816_/B _5945_/Y vssd1 vssd1 vccd1 vccd1 _6044_/Y sky130_fd_sc_hd__a21oi_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3256_/A vssd1 vssd1 vccd1 vccd1 _4540_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_85_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3187_ input8/X vssd1 vssd1 vccd1 vccd1 _3441_/A sky130_fd_sc_hd__inv_2
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5828_ _5816_/B _5802_/A _5944_/A vssd1 vssd1 vccd1 vccd1 _5828_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5759_ _5672_/X _5685_/X _5786_/A _5786_/B vssd1 vssd1 vccd1 vccd1 _5759_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_89_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4090_ _4090_/A _4625_/A _4890_/C vssd1 vssd1 vccd1 vccd1 _4091_/B sky130_fd_sc_hd__nand3_2
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4992_ _4549_/X _4689_/X _4720_/Y _4975_/B vssd1 vssd1 vccd1 vccd1 _5004_/B sky130_fd_sc_hd__o31a_2
X_3943_ _3780_/X _3778_/A _3819_/B vssd1 vssd1 vccd1 vccd1 _3943_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3874_ _3868_/Y _3872_/Y _3873_/Y vssd1 vssd1 vccd1 vccd1 _3875_/C sky130_fd_sc_hd__a21o_1
X_5613_ _5267_/B _5268_/A _5370_/X vssd1 vssd1 vccd1 vccd1 _5613_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_31_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5544_ _4287_/B _5453_/B _5554_/A vssd1 vssd1 vccd1 vccd1 _5549_/A sky130_fd_sc_hd__o21ai_1
X_5475_ _5475_/A _5475_/B vssd1 vssd1 vccd1 vccd1 _5479_/B sky130_fd_sc_hd__nor2_1
X_4426_ _4489_/A _4489_/B vssd1 vssd1 vccd1 vccd1 _4468_/A sky130_fd_sc_hd__nand2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ input6/X vssd1 vssd1 vccd1 vccd1 _4387_/A sky130_fd_sc_hd__inv_2
X_4288_ _4285_/Y _4287_/Y _4284_/C vssd1 vssd1 vccd1 vccd1 _4288_/Y sky130_fd_sc_hd__a21oi_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ _3300_/C _3300_/D _3306_/Y vssd1 vssd1 vccd1 vccd1 _3309_/C sky130_fd_sc_hd__a21o_1
XFILLER_86_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6027_ _6021_/A _6110_/B vssd1 vssd1 vccd1 vccd1 _6027_/X sky130_fd_sc_hd__and2b_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _3240_/A _3240_/B _3240_/C vssd1 vssd1 vccd1 vccd1 _3241_/A sky130_fd_sc_hd__a21o_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3590_ _3597_/B vssd1 vssd1 vccd1 vccd1 _3857_/C sky130_fd_sc_hd__inv_2
X_5260_ _5051_/Y _5259_/X _5056_/C _5082_/A vssd1 vssd1 vccd1 vccd1 _5260_/Y sky130_fd_sc_hd__a2bb2oi_2
X_4211_ _4211_/A _4211_/B vssd1 vssd1 vccd1 vccd1 _4220_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5191_ _5012_/B _5012_/C _5012_/A vssd1 vssd1 vccd1 vccd1 _5191_/Y sky130_fd_sc_hd__a21oi_1
X_4142_ _4054_/A _4054_/B _4054_/C vssd1 vssd1 vccd1 vccd1 _4142_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4073_ _4571_/A _4571_/B _5212_/B _5541_/B vssd1 vssd1 vccd1 vccd1 _4073_/Y sky130_fd_sc_hd__nand4_4
XFILLER_36_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4975_ _4975_/A _4975_/B _4975_/C vssd1 vssd1 vccd1 vccd1 _4976_/B sky130_fd_sc_hd__nand3_1
X_3926_ _3927_/A _4128_/B _3927_/C vssd1 vssd1 vccd1 vccd1 _3928_/B sky130_fd_sc_hd__a21o_1
X_3857_ _3857_/A _3857_/B _3857_/C vssd1 vssd1 vccd1 vccd1 _3857_/X sky130_fd_sc_hd__and3_1
X_3788_ _5029_/A vssd1 vssd1 vccd1 vccd1 _4904_/B sky130_fd_sc_hd__buf_2
X_5527_ _5527_/A vssd1 vssd1 vccd1 vccd1 _5629_/A sky130_fd_sc_hd__inv_2
X_5458_ _5460_/A _5460_/B _5468_/C _5468_/D vssd1 vssd1 vccd1 vccd1 _5458_/Y sky130_fd_sc_hd__nand4_2
X_4409_ _4088_/Y _4257_/Y _4406_/Y _4408_/Y vssd1 vssd1 vccd1 vccd1 _4409_/X sky130_fd_sc_hd__o22a_1
X_5389_ _5246_/X _5379_/A _5375_/Y vssd1 vssd1 vccd1 vccd1 _5391_/A sky130_fd_sc_hd__o21ai_1
XFILLER_75_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4760_ _4574_/Y _4577_/Y _4598_/A _4587_/A vssd1 vssd1 vccd1 vccd1 _4765_/B sky130_fd_sc_hd__a2bb2oi_4
X_3711_ _3711_/A vssd1 vssd1 vccd1 vccd1 _4936_/A sky130_fd_sc_hd__clkbuf_4
X_4691_ _3543_/B _4530_/C _5701_/A _4700_/A vssd1 vssd1 vccd1 vccd1 _4691_/Y sky130_fd_sc_hd__a22oi_2
X_3642_ _3639_/X _3641_/X _3691_/A _3625_/Y vssd1 vssd1 vccd1 vccd1 _3720_/B sky130_fd_sc_hd__o211ai_2
X_5312_ _5289_/Y _5293_/Y _5297_/Y _5304_/B vssd1 vssd1 vccd1 vccd1 _5313_/C sky130_fd_sc_hd__o211ai_1
X_3573_ _3736_/A _3736_/B _3736_/C vssd1 vssd1 vccd1 vccd1 _3607_/B sky130_fd_sc_hd__nand3_2
X_6292_ _6283_/X _6292_/B _6292_/C vssd1 vssd1 vccd1 vccd1 _6292_/Y sky130_fd_sc_hd__nand3b_4
X_5243_ _5268_/A _5268_/B vssd1 vssd1 vccd1 vccd1 _5420_/A sky130_fd_sc_hd__nand2_1
X_5174_ _5004_/B _5021_/B _4991_/Y vssd1 vssd1 vccd1 vccd1 _5180_/A sky130_fd_sc_hd__a21oi_2
X_4125_ _4133_/A _4133_/B _4141_/A vssd1 vssd1 vccd1 vccd1 _4125_/Y sky130_fd_sc_hd__nand3_2
XFILLER_56_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4056_ _4852_/A _4590_/B vssd1 vssd1 vccd1 vccd1 _4071_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4958_ _4958_/A _4958_/B _5532_/C _5299_/D vssd1 vssd1 vccd1 vccd1 _4958_/X sky130_fd_sc_hd__and4_2
XFILLER_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3909_ _3747_/B _3889_/A _4868_/A _5123_/A _3891_/Y vssd1 vssd1 vccd1 vccd1 _3911_/B
+ sky130_fd_sc_hd__o2111ai_1
X_4889_ _5448_/B vssd1 vssd1 vccd1 vccd1 _5810_/A sky130_fd_sc_hd__buf_4
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5930_ _5407_/C _6016_/A _5986_/B _5809_/A vssd1 vssd1 vccd1 vccd1 _5933_/A sky130_fd_sc_hd__a22o_1
XFILLER_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5861_ _5822_/Y _5944_/B _5827_/Y _5828_/X vssd1 vssd1 vccd1 vccd1 _5865_/A sky130_fd_sc_hd__o211ai_1
XFILLER_33_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5792_ _5792_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _5793_/B sky130_fd_sc_hd__nand2_1
X_4812_ _4660_/B _4645_/Y _4639_/Y vssd1 vssd1 vccd1 vccd1 _4815_/A sky130_fd_sc_hd__a21boi_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4743_ _4568_/A _4568_/B _4576_/A vssd1 vssd1 vccd1 vccd1 _4743_/X sky130_fd_sc_hd__o21a_1
X_4674_ _6235_/A vssd1 vssd1 vccd1 vccd1 _4674_/X sky130_fd_sc_hd__clkbuf_4
X_3625_ _3625_/A _3625_/B _3625_/C vssd1 vssd1 vccd1 vccd1 _3625_/Y sky130_fd_sc_hd__nand3_4
X_3556_ _3552_/Y _3554_/Y _3555_/Y vssd1 vssd1 vccd1 vccd1 _3559_/B sky130_fd_sc_hd__a21o_1
X_6275_ _6277_/A _6275_/B _6275_/C vssd1 vssd1 vccd1 vccd1 _6275_/Y sky130_fd_sc_hd__nor3_1
X_5226_ _5281_/A _5271_/A _5281_/C vssd1 vssd1 vccd1 vccd1 _5226_/X sky130_fd_sc_hd__and3_1
X_3487_ _3487_/A vssd1 vssd1 vccd1 vccd1 _3592_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5157_ _5325_/A _5157_/B _5200_/A _5200_/B vssd1 vssd1 vccd1 vccd1 _5159_/B sky130_fd_sc_hd__nand4_1
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4108_ _4700_/A vssd1 vssd1 vccd1 vccd1 _5302_/C sky130_fd_sc_hd__clkbuf_4
X_5088_ _5088_/A _5088_/B vssd1 vssd1 vccd1 vccd1 _5088_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4039_ _4029_/Y _4032_/Y _3964_/B _4036_/Y _4038_/Y vssd1 vssd1 vccd1 vccd1 _4041_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_72_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4390_ _4390_/A _5302_/B vssd1 vssd1 vccd1 vccd1 _4390_/Y sky130_fd_sc_hd__nand2_2
X_3410_ _3410_/A _3410_/B vssd1 vssd1 vccd1 vccd1 _3486_/C sky130_fd_sc_hd__xnor2_2
X_3341_ _4432_/A _3542_/A vssd1 vssd1 vccd1 vccd1 _3342_/B sky130_fd_sc_hd__nand2_4
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6060_/A _6193_/B vssd1 vssd1 vccd1 vccd1 _6060_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3272_ _5053_/A _3356_/A vssd1 vssd1 vccd1 vccd1 _3276_/A sky130_fd_sc_hd__nand2_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _4711_/B _5010_/X _5001_/Y _5005_/Y vssd1 vssd1 vccd1 vccd1 _5012_/C sky130_fd_sc_hd__o211ai_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5913_ _5914_/A _5914_/B _5914_/C _5998_/B vssd1 vssd1 vccd1 vccd1 _5989_/A sky130_fd_sc_hd__a22o_1
XFILLER_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5844_ _6124_/B vssd1 vssd1 vccd1 vccd1 _6203_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_21_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5775_ _5974_/A _5974_/B vssd1 vssd1 vccd1 vccd1 _5780_/A sky130_fd_sc_hd__nand2_1
X_4726_ _4721_/X _4722_/Y _4719_/Y _4712_/Y vssd1 vssd1 vccd1 vccd1 _4975_/B sky130_fd_sc_hd__o211ai_2
X_4657_ _4659_/A _4659_/B _4649_/Y _4650_/Y _4645_/Y vssd1 vssd1 vccd1 vccd1 _4661_/B
+ sky130_fd_sc_hd__o221ai_4
X_3608_ _3574_/A _3574_/C _3574_/B _3486_/B _3479_/A vssd1 vssd1 vccd1 vccd1 _3609_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4588_ _4574_/Y _4577_/Y _4606_/C vssd1 vssd1 vccd1 vccd1 _4599_/A sky130_fd_sc_hd__o21ai_1
XFILLER_88_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3539_ _3525_/Y _3526_/X _3535_/Y _3538_/X vssd1 vssd1 vccd1 vccd1 _3540_/A sky130_fd_sc_hd__o211ai_2
XFILLER_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6258_ _6258_/A _6258_/B _6258_/C vssd1 vssd1 vccd1 vccd1 _6258_/X sky130_fd_sc_hd__or3_1
XFILLER_88_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6189_ _6190_/C _6214_/A _6190_/A vssd1 vssd1 vccd1 vccd1 _6224_/A sky130_fd_sc_hd__o21a_1
XFILLER_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5209_ _5209_/A _5575_/A _5541_/B _5211_/B vssd1 vssd1 vccd1 vccd1 _5209_/Y sky130_fd_sc_hd__nand4_2
XFILLER_29_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3890_ _4730_/A _4906_/B vssd1 vssd1 vccd1 vccd1 _4064_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5560_ _5694_/A _5694_/B _5561_/C _5694_/C vssd1 vssd1 vccd1 vccd1 _5563_/A sky130_fd_sc_hd__a22o_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5491_ _5634_/B _5480_/Y _5477_/A _5623_/B _5624_/A vssd1 vssd1 vccd1 vccd1 _5493_/B
+ sky130_fd_sc_hd__o2111ai_1
X_4511_ _4511_/A _4511_/B _4506_/B vssd1 vssd1 vccd1 vccd1 _4511_/Y sky130_fd_sc_hd__nor3b_1
X_4442_ _4057_/X _4429_/A _4435_/Y vssd1 vssd1 vccd1 vccd1 _4442_/X sky130_fd_sc_hd__o21a_1
X_4373_ _5446_/A vssd1 vssd1 vccd1 vccd1 _5453_/B sky130_fd_sc_hd__clkbuf_4
X_6112_ _6112_/A _6112_/B _6112_/C vssd1 vssd1 vccd1 vccd1 _6219_/C sky130_fd_sc_hd__nand3_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _5064_/A vssd1 vssd1 vccd1 vccd1 _5248_/A sky130_fd_sc_hd__buf_4
X_6043_ _5942_/C _5942_/B _5942_/A _5940_/C vssd1 vssd1 vccd1 vccd1 _6043_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _4193_/A _3960_/B _3677_/A _5372_/B vssd1 vssd1 vccd1 vccd1 _3265_/D sky130_fd_sc_hd__nand4_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _3186_/A vssd1 vssd1 vccd1 vccd1 _3186_/X sky130_fd_sc_hd__buf_2
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5827_ _5673_/B _5690_/X _5825_/X _5826_/Y vssd1 vssd1 vccd1 vccd1 _5827_/Y sky130_fd_sc_hd__o2bb2ai_2
X_5758_ _5625_/A _5625_/B _5625_/D _5619_/Y vssd1 vssd1 vccd1 vccd1 _5761_/B sky130_fd_sc_hd__a31oi_4
X_4709_ _4547_/A _4708_/C _5532_/D _4540_/B vssd1 vssd1 vccd1 vccd1 _4711_/B sky130_fd_sc_hd__a22oi_4
X_5689_ _5834_/A vssd1 vssd1 vccd1 vccd1 _5852_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4991_ _4990_/Y _4985_/Y _4979_/Y vssd1 vssd1 vccd1 vccd1 _4991_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_16_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3942_ _3752_/X _3757_/X _3809_/B _3809_/A vssd1 vssd1 vccd1 vccd1 _3942_/X sky130_fd_sc_hd__o211a_1
XFILLER_31_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3873_ _4708_/A _4779_/B vssd1 vssd1 vccd1 vccd1 _3873_/Y sky130_fd_sc_hd__nand2_2
X_5612_ _5612_/A _5612_/B vssd1 vssd1 vccd1 vccd1 _5612_/X sky130_fd_sc_hd__and2_1
X_5543_ _5538_/X _5540_/X _5542_/Y vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__o21ai_1
X_5474_ _5479_/A _5634_/A _5475_/B _5475_/A vssd1 vssd1 vccd1 vccd1 _5477_/A sky130_fd_sc_hd__o2bb2ai_1
X_4425_ _4414_/X _4420_/X _4422_/X _4424_/X vssd1 vssd1 vccd1 vccd1 _4489_/B sky130_fd_sc_hd__o2bb2ai_1
X_4356_ _4356_/A vssd1 vssd1 vccd1 vccd1 _4362_/B sky130_fd_sc_hd__clkbuf_2
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ _3304_/Y _3305_/Y _3300_/C _3306_/Y vssd1 vssd1 vccd1 vccd1 _3309_/B sky130_fd_sc_hd__o211ai_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _5603_/A _4287_/B vssd1 vssd1 vccd1 vccd1 _4287_/Y sky130_fd_sc_hd__nor2_2
X_6026_ _6025_/X _5942_/A _5942_/B vssd1 vssd1 vccd1 vccd1 _6037_/B sky130_fd_sc_hd__o21a_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3238_ _3199_/C _3236_/Y _3237_/X vssd1 vssd1 vccd1 vccd1 _3240_/C sky130_fd_sc_hd__o21a_1
XFILLER_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3169_ _3165_/X _3167_/Y _3310_/A _3229_/D vssd1 vssd1 vccd1 vccd1 _3170_/B sky130_fd_sc_hd__o211a_2
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4210_ _4194_/Y _4198_/Y _4219_/B vssd1 vssd1 vccd1 vccd1 _4210_/Y sky130_fd_sc_hd__o21ai_1
X_5190_ _5190_/A _5190_/B vssd1 vssd1 vccd1 vccd1 _5190_/Y sky130_fd_sc_hd__nor2_1
X_4141_ _4141_/A _4141_/B _4141_/C vssd1 vssd1 vccd1 vccd1 _4141_/Y sky130_fd_sc_hd__nand3_1
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4072_ _4590_/B vssd1 vssd1 vccd1 vccd1 _5541_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4974_ _4549_/X _4689_/X _4720_/Y _4723_/X vssd1 vssd1 vccd1 vccd1 _4976_/A sky130_fd_sc_hd__o22ai_1
X_3925_ _3918_/C _3923_/Y _3924_/Y vssd1 vssd1 vccd1 vccd1 _3927_/C sky130_fd_sc_hd__a21oi_2
X_3856_ _3856_/A _3856_/B vssd1 vssd1 vccd1 vccd1 _3856_/Y sky130_fd_sc_hd__nor2_1
X_3787_ _3787_/A _3787_/B vssd1 vssd1 vccd1 vccd1 _3791_/A sky130_fd_sc_hd__nand2_1
X_5526_ _5479_/A _5479_/B _5480_/Y vssd1 vssd1 vccd1 vccd1 _5527_/A sky130_fd_sc_hd__a21oi_1
X_5457_ _5457_/A _5457_/B _5457_/C vssd1 vssd1 vccd1 vccd1 _5468_/D sky130_fd_sc_hd__nand3_2
X_4408_ _5378_/A _4777_/C _5284_/C _3551_/A vssd1 vssd1 vccd1 vccd1 _4408_/Y sky130_fd_sc_hd__a22oi_2
X_5388_ _5390_/A _6202_/B _5246_/X _5598_/A _5375_/Y vssd1 vssd1 vccd1 vccd1 _5388_/Y
+ sky130_fd_sc_hd__o221ai_4
X_4339_ _4163_/B _3998_/D _4163_/Y _3859_/B vssd1 vssd1 vccd1 vccd1 _4339_/X sky130_fd_sc_hd__o22a_1
XFILLER_86_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6009_ _6009_/A vssd1 vssd1 vccd1 vccd1 _6127_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3710_ _3350_/Y _5867_/A _3611_/X _3679_/Y _3676_/Y vssd1 vssd1 vccd1 vccd1 _3710_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4690_ _4958_/A _5704_/B vssd1 vssd1 vccd1 vccd1 _4690_/Y sky130_fd_sc_hd__nand2_1
X_3641_ _3641_/A _4422_/B _4362_/C vssd1 vssd1 vccd1 vccd1 _3641_/X sky130_fd_sc_hd__and3_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3572_ _3576_/A _3730_/B _3577_/B _3703_/B vssd1 vssd1 vccd1 vccd1 _3736_/C sky130_fd_sc_hd__nand4_2
X_5311_ _5303_/A _5303_/B _5304_/A vssd1 vssd1 vccd1 vccd1 _5313_/B sky130_fd_sc_hd__o21ai_1
X_6291_ _6289_/B _6289_/C _6289_/A vssd1 vssd1 vccd1 vccd1 _6292_/C sky130_fd_sc_hd__a21o_1
X_5242_ _5258_/A _5046_/B _5239_/Y _5240_/X _5241_/X vssd1 vssd1 vccd1 vccd1 _5268_/B
+ sky130_fd_sc_hd__o221ai_4
X_5173_ _5173_/A vssd1 vssd1 vccd1 vccd1 _5182_/A sky130_fd_sc_hd__clkbuf_2
X_4124_ _4124_/A _4124_/B _4124_/C vssd1 vssd1 vccd1 vccd1 _4141_/A sky130_fd_sc_hd__nand3_2
XFILLER_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput1 a[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
XFILLER_28_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4055_ _4078_/A vssd1 vssd1 vccd1 vccd1 _4590_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_64_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4957_ _4939_/A _5302_/C _5810_/B _5805_/B _4956_/X vssd1 vssd1 vccd1 vccd1 _4957_/X
+ sky130_fd_sc_hd__a41o_2
X_3908_ _3908_/A vssd1 vssd1 vccd1 vccd1 _4868_/A sky130_fd_sc_hd__buf_2
X_4888_ _4752_/A _4754_/A _4758_/C vssd1 vssd1 vccd1 vccd1 _4891_/A sky130_fd_sc_hd__a21o_1
X_3839_ _3833_/X _3839_/B _3839_/C vssd1 vssd1 vccd1 vccd1 _3847_/C sky130_fd_sc_hd__nand3b_1
XFILLER_20_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5509_ _5509_/A _5514_/C _5509_/C vssd1 vssd1 vccd1 vccd1 _5643_/B sky130_fd_sc_hd__nand3_1
XFILLER_10_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5860_ _5860_/A _5860_/B _5860_/C vssd1 vssd1 vccd1 vccd1 _5860_/Y sky130_fd_sc_hd__nand3_1
XFILLER_80_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4811_ _4996_/A _4996_/B _4995_/A vssd1 vssd1 vccd1 vccd1 _4822_/B sky130_fd_sc_hd__nand3_2
X_5791_ _5704_/Y _5706_/Y _5698_/Y vssd1 vssd1 vccd1 vccd1 _5791_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4742_ _4742_/A vssd1 vssd1 vccd1 vccd1 _4742_/X sky130_fd_sc_hd__clkbuf_2
X_4673_ _6171_/C vssd1 vssd1 vccd1 vccd1 _6235_/A sky130_fd_sc_hd__clkbuf_4
X_3624_ _3617_/A _3630_/B _3623_/Y vssd1 vssd1 vccd1 vccd1 _3625_/C sky130_fd_sc_hd__a21o_1
X_3555_ _3555_/A _4236_/A vssd1 vssd1 vccd1 vccd1 _3555_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6274_ _6274_/A vssd1 vssd1 vccd1 vccd1 _6274_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3486_ _3486_/A _3486_/B _3486_/C vssd1 vssd1 vccd1 vccd1 _3584_/B sky130_fd_sc_hd__nand3_1
X_5225_ _5224_/Y _5026_/Y _5220_/Y vssd1 vssd1 vccd1 vccd1 _5281_/C sky130_fd_sc_hd__a21oi_2
X_5156_ _4965_/X _5152_/X _5149_/A _5145_/A vssd1 vssd1 vccd1 vccd1 _5200_/B sky130_fd_sc_hd__o211ai_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4107_ _3898_/X _3923_/Y _4105_/Y _4106_/X vssd1 vssd1 vccd1 vccd1 _4135_/C sky130_fd_sc_hd__o211ai_4
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5087_ _5087_/A _5087_/B _5087_/C _5919_/B vssd1 vssd1 vccd1 vccd1 _5087_/X sky130_fd_sc_hd__and4_1
X_4038_ _4038_/A _4038_/B _4201_/A vssd1 vssd1 vccd1 vccd1 _4038_/Y sky130_fd_sc_hd__nand3_1
XFILLER_64_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _5989_/A _6024_/A vssd1 vssd1 vccd1 vccd1 _5989_/Y sky130_fd_sc_hd__nand2_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3340_ _3348_/B vssd1 vssd1 vccd1 vccd1 _3358_/D sky130_fd_sc_hd__clkbuf_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _4711_/A _6235_/A _5006_/Y _5007_/Y vssd1 vssd1 vccd1 vccd1 _5010_/X sky130_fd_sc_hd__o22a_1
X_3271_ _4738_/A vssd1 vssd1 vccd1 vccd1 _5053_/A sky130_fd_sc_hd__clkbuf_4
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5912_ _5912_/A _5912_/B vssd1 vssd1 vccd1 vccd1 _5949_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5843_ _5994_/A _6065_/C _6065_/D _5905_/A vssd1 vssd1 vccd1 vccd1 _5843_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5774_ _5773_/B _5773_/C _5773_/A vssd1 vssd1 vccd1 vccd1 _5974_/B sky130_fd_sc_hd__a21o_1
X_4725_ _4712_/Y _4988_/B _4719_/Y vssd1 vssd1 vccd1 vccd1 _4975_/A sky130_fd_sc_hd__a21o_1
X_4656_ _4564_/X _4561_/X _4554_/Y _4560_/A vssd1 vssd1 vccd1 vccd1 _4659_/B sky130_fd_sc_hd__o211a_1
X_3607_ _3607_/A _3607_/B _3607_/C vssd1 vssd1 vccd1 vccd1 _3607_/Y sky130_fd_sc_hd__nand3_1
X_4587_ _4587_/A vssd1 vssd1 vccd1 vccd1 _4606_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3538_ _3658_/A _3657_/B _3657_/A vssd1 vssd1 vccd1 vccd1 _3538_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6257_ _6257_/A _6257_/B _6257_/C vssd1 vssd1 vccd1 vccd1 _6258_/C sky130_fd_sc_hd__and3_1
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3469_ _4711_/A _5390_/A _3368_/B _3552_/A _3419_/Y vssd1 vssd1 vccd1 vccd1 _3471_/A
+ sky130_fd_sc_hd__o221a_1
X_6188_ _6156_/A _6156_/B _6156_/C vssd1 vssd1 vccd1 vccd1 _6190_/A sky130_fd_sc_hd__a21boi_2
X_5208_ _5208_/A _5208_/B vssd1 vssd1 vccd1 vccd1 _5208_/Y sky130_fd_sc_hd__nand2_4
X_5139_ _5126_/Y _5366_/A _5138_/Y vssd1 vssd1 vccd1 vccd1 _5139_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_72_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5490_ _5490_/A _5490_/B _5490_/C _5490_/D vssd1 vssd1 vccd1 vccd1 _5623_/B sky130_fd_sc_hd__nand4_1
X_4510_ _4333_/A _4333_/C _4333_/B vssd1 vssd1 vccd1 vccd1 _4511_/B sky130_fd_sc_hd__a21boi_1
XFILLER_7_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4441_ _4601_/A _4601_/B _4441_/C vssd1 vssd1 vccd1 vccd1 _4463_/A sky130_fd_sc_hd__nand3_4
X_6111_ _5933_/B _5987_/Y _6051_/B _6049_/B _6049_/A vssd1 vssd1 vccd1 vccd1 _6112_/C
+ sky130_fd_sc_hd__a32o_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4372_ _4372_/A vssd1 vssd1 vccd1 vccd1 _5446_/A sky130_fd_sc_hd__clkbuf_4
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _4884_/A vssd1 vssd1 vccd1 vccd1 _5064_/A sky130_fd_sc_hd__buf_2
X_6042_ _5860_/C _5989_/Y _5960_/B _6041_/Y vssd1 vssd1 vccd1 vccd1 _6047_/B sky130_fd_sc_hd__o211ai_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _3414_/B vssd1 vssd1 vccd1 vccd1 _5372_/B sky130_fd_sc_hd__clkbuf_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3185_ _4176_/A vssd1 vssd1 vccd1 vccd1 _3186_/A sky130_fd_sc_hd__inv_2
XFILLER_26_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5826_ _5826_/A _5826_/B vssd1 vssd1 vccd1 vccd1 _5826_/Y sky130_fd_sc_hd__nand2_1
X_5757_ _5693_/X _5747_/Y _5756_/Y vssd1 vssd1 vccd1 vccd1 _5761_/A sky130_fd_sc_hd__o21ai_1
X_4708_ _4708_/A _4708_/B _4708_/C _5299_/D vssd1 vssd1 vccd1 vccd1 _4711_/D sky130_fd_sc_hd__and4_2
X_5688_ _5688_/A vssd1 vssd1 vccd1 vccd1 _6137_/C sky130_fd_sc_hd__clkbuf_2
X_4639_ _4639_/A _4639_/B _4639_/C vssd1 vssd1 vccd1 vccd1 _4639_/Y sky130_fd_sc_hd__nand3_1
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4990_ _4980_/Y _4982_/Y _4972_/Y _4989_/Y vssd1 vssd1 vccd1 vccd1 _4990_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3941_ _3938_/A _3938_/B _3939_/A vssd1 vssd1 vccd1 vccd1 _4008_/A sky130_fd_sc_hd__o21ai_1
XFILLER_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3872_ _4708_/B _4700_/A _4788_/A _4238_/D vssd1 vssd1 vccd1 vccd1 _3872_/Y sky130_fd_sc_hd__nand4_4
X_5611_ _5611_/A _5611_/B vssd1 vssd1 vccd1 vccd1 _5616_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5542_ _5542_/A _5542_/B vssd1 vssd1 vccd1 vccd1 _5542_/Y sky130_fd_sc_hd__nand2_2
XFILLER_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5473_ _5297_/B _5297_/C _5297_/A vssd1 vssd1 vccd1 vccd1 _5475_/A sky130_fd_sc_hd__a21oi_2
X_4424_ _5347_/A _5831_/A _5435_/A _5669_/A vssd1 vssd1 vccd1 vccd1 _4424_/X sky130_fd_sc_hd__and4_1
X_4355_ _4355_/A _4355_/B _4708_/C _5299_/D vssd1 vssd1 vccd1 vccd1 _4356_/A sky130_fd_sc_hd__nand4_2
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ _3306_/A _3306_/B vssd1 vssd1 vccd1 vccd1 _3306_/Y sky130_fd_sc_hd__nand2_1
X_4286_ _5034_/B vssd1 vssd1 vccd1 vccd1 _4287_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_58_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6025_ _6025_/A _6025_/B _6025_/C vssd1 vssd1 vccd1 vccd1 _6025_/X sky130_fd_sc_hd__and3_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _3966_/B _3310_/C _5845_/A _3521_/A vssd1 vssd1 vccd1 vccd1 _3237_/X sky130_fd_sc_hd__a22o_1
X_3168_ _3310_/A _3229_/D _3165_/X _3167_/Y vssd1 vssd1 vccd1 vccd1 _3170_/A sky130_fd_sc_hd__a211oi_4
XFILLER_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5809_ _5809_/A _5809_/B vssd1 vssd1 vccd1 vccd1 _5809_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4140_ _3984_/A _3984_/C _3945_/A vssd1 vssd1 vccd1 vccd1 _4141_/C sky130_fd_sc_hd__a21boi_1
X_4071_ _4071_/A _4071_/B vssd1 vssd1 vccd1 vccd1 _4071_/Y sky130_fd_sc_hd__nand2_2
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4973_ _4984_/A _4984_/B _4972_/Y vssd1 vssd1 vccd1 vccd1 _4973_/Y sky130_fd_sc_hd__o21ai_2
X_3924_ _4236_/A _5299_/A _3918_/B _3918_/C vssd1 vssd1 vccd1 vccd1 _3924_/Y sky130_fd_sc_hd__a22oi_1
X_3855_ _4163_/A _4163_/B vssd1 vssd1 vccd1 vccd1 _3859_/A sky130_fd_sc_hd__nand2_1
X_3786_ _4184_/A _5209_/A vssd1 vssd1 vccd1 vccd1 _3787_/B sky130_fd_sc_hd__nand2_2
X_5525_ _5525_/A _5525_/B vssd1 vssd1 vccd1 vccd1 _5631_/A sky130_fd_sc_hd__nand2_1
X_5456_ _5453_/A _6236_/A _5291_/X _5542_/A _5445_/Y vssd1 vssd1 vccd1 vccd1 _5457_/C
+ sky130_fd_sc_hd__o221ai_2
XFILLER_59_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4407_ _4407_/A vssd1 vssd1 vccd1 vccd1 _4777_/C sky130_fd_sc_hd__clkbuf_2
X_5387_ _3179_/C _5676_/A _4747_/A vssd1 vssd1 vccd1 vccd1 _5387_/X sky130_fd_sc_hd__a21o_1
X_4338_ _4338_/A _4520_/B vssd1 vssd1 vccd1 vccd1 _4338_/Y sky130_fd_sc_hd__nand2_1
X_4269_ _4901_/B vssd1 vssd1 vccd1 vccd1 _4761_/B sky130_fd_sc_hd__buf_2
X_6008_ _6005_/Y _6006_/X _6007_/X vssd1 vssd1 vccd1 vccd1 _6091_/A sky130_fd_sc_hd__o21bai_4
XFILLER_82_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3640_ _4390_/A vssd1 vssd1 vccd1 vccd1 _4362_/C sky130_fd_sc_hd__buf_2
X_3571_ _3478_/A _3570_/Y _3486_/A _3486_/C vssd1 vssd1 vccd1 vccd1 _3736_/B sky130_fd_sc_hd__a22o_1
X_6290_ _6290_/A _6290_/B vssd1 vssd1 vccd1 vccd1 _6290_/Y sky130_fd_sc_hd__nor2_1
X_5310_ _5310_/A _5310_/B vssd1 vssd1 vccd1 vccd1 _5313_/A sky130_fd_sc_hd__nand2_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5241_ _5258_/A _5046_/B _5060_/Y vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__a21o_1
X_5172_ _5172_/A _5172_/B _5172_/C vssd1 vssd1 vccd1 vccd1 _5173_/A sky130_fd_sc_hd__nand3_2
XFILLER_68_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4123_ _4124_/C _4124_/A _4124_/B vssd1 vssd1 vccd1 vccd1 _4123_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_83_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput2 a[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_4
X_4054_ _4054_/A _4054_/B _4054_/C vssd1 vssd1 vccd1 vccd1 _4054_/X sky130_fd_sc_hd__and3_2
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4956_ _4956_/A _5134_/B vssd1 vssd1 vccd1 vccd1 _4956_/X sky130_fd_sc_hd__and2_2
X_3907_ _3441_/A _4460_/B _3895_/A vssd1 vssd1 vccd1 vccd1 _3911_/A sky130_fd_sc_hd__o21ai_1
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4887_ _4885_/X _4886_/Y _4865_/Y _4871_/X vssd1 vssd1 vccd1 vccd1 _4893_/B sky130_fd_sc_hd__o211ai_1
X_3838_ _3837_/C _3837_/A _3837_/B vssd1 vssd1 vccd1 vccd1 _3839_/C sky130_fd_sc_hd__a21o_1
X_5508_ _5514_/C _5643_/A _5509_/A vssd1 vssd1 vccd1 vccd1 _5510_/C sky130_fd_sc_hd__a21o_1
X_3769_ _3897_/A vssd1 vssd1 vccd1 vccd1 _5378_/A sky130_fd_sc_hd__buf_4
X_5439_ _5465_/C _4829_/A _5438_/Y vssd1 vssd1 vccd1 vccd1 _5460_/A sky130_fd_sc_hd__a21o_1
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _4793_/X _4798_/Y _4803_/Y _4814_/B vssd1 vssd1 vccd1 vccd1 _4995_/A sky130_fd_sc_hd__o211ai_2
X_5790_ _6125_/A _6124_/A _5688_/A _6010_/B _5789_/Y vssd1 vssd1 vccd1 vccd1 _5790_/X
+ sky130_fd_sc_hd__a41o_1
X_4741_ _4741_/A _4741_/B _4741_/C vssd1 vssd1 vccd1 vccd1 _4742_/A sky130_fd_sc_hd__nand3_1
X_4672_ _4390_/Y _4386_/Y _4362_/B _4680_/C _4680_/D vssd1 vssd1 vccd1 vccd1 _4672_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_3623_ _4542_/A _5401_/A vssd1 vssd1 vccd1 vccd1 _3623_/Y sky130_fd_sc_hd__nand2_1
X_3554_ _5251_/A _4708_/B _5373_/A _4958_/B vssd1 vssd1 vccd1 vccd1 _3554_/Y sky130_fd_sc_hd__nand4_2
X_6273_ _6273_/A _6273_/B vssd1 vssd1 vccd1 vccd1 _6273_/Y sky130_fd_sc_hd__nand2_4
X_3485_ _3486_/A _3486_/B _3486_/C vssd1 vssd1 vccd1 vccd1 _3584_/A sky130_fd_sc_hd__a21o_1
XFILLER_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5224_ _5834_/A _5808_/A vssd1 vssd1 vccd1 vccd1 _5224_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5155_ _5145_/A _5149_/A _5150_/Y vssd1 vssd1 vccd1 vccd1 _5200_/A sky130_fd_sc_hd__a21o_1
XFILLER_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5086_ _5570_/A vssd1 vssd1 vccd1 vccd1 _5919_/B sky130_fd_sc_hd__buf_2
X_4106_ _5134_/A _3795_/B _4302_/A _4105_/B vssd1 vssd1 vccd1 vccd1 _4106_/X sky130_fd_sc_hd__a22o_1
XFILLER_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4037_ _4020_/A _4020_/B _4182_/A _4025_/Y vssd1 vssd1 vccd1 vccd1 _4038_/A sky130_fd_sc_hd__o2bb2ai_1
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5988_ _5957_/A _5957_/B _5957_/C _5961_/X vssd1 vssd1 vccd1 vccd1 _6049_/A sky130_fd_sc_hd__a31o_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4939_ _4939_/A _5302_/C _5810_/B _5809_/B vssd1 vssd1 vccd1 vccd1 _4943_/B sky130_fd_sc_hd__nand4_2
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _4067_/A _3270_/B _4547_/A _4958_/B vssd1 vssd1 vccd1 vccd1 _3345_/B sky130_fd_sc_hd__nand4_4
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5911_ _5911_/A _5911_/B vssd1 vssd1 vccd1 vccd1 _5912_/B sky130_fd_sc_hd__nor2_1
XFILLER_34_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5842_ _5842_/A vssd1 vssd1 vccd1 vccd1 _6065_/C sky130_fd_sc_hd__clkbuf_2
X_5773_ _5773_/A _5773_/B _5773_/C vssd1 vssd1 vccd1 vccd1 _5974_/A sky130_fd_sc_hd__nand3_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4724_ _4549_/X _4689_/X _4720_/Y _4723_/X vssd1 vssd1 vccd1 vccd1 _4809_/A sky130_fd_sc_hd__o22a_1
X_4655_ _4554_/Y _4817_/A _4562_/X vssd1 vssd1 vccd1 vccd1 _4659_/A sky130_fd_sc_hd__a21oi_2
X_3606_ _3593_/B _3488_/X _3605_/Y vssd1 vssd1 vccd1 vccd1 _3606_/Y sky130_fd_sc_hd__a21oi_1
X_4586_ _4586_/A _4586_/B _4586_/C vssd1 vssd1 vccd1 vccd1 _4587_/A sky130_fd_sc_hd__nand3_1
X_3537_ _5229_/A _4532_/A vssd1 vssd1 vccd1 vccd1 _3657_/A sky130_fd_sc_hd__nand2_1
X_6256_ _6260_/A _6260_/B vssd1 vssd1 vccd1 vccd1 _6258_/B sky130_fd_sc_hd__nor2_1
X_3468_ _3468_/A vssd1 vssd1 vccd1 vccd1 _4711_/A sky130_fd_sc_hd__buf_2
X_6187_ _6187_/A _6222_/A _6187_/C vssd1 vssd1 vccd1 vccd1 _6214_/A sky130_fd_sc_hd__nor3_2
X_3399_ _4901_/A vssd1 vssd1 vccd1 vccd1 _5397_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5207_ _5207_/A _5207_/B vssd1 vssd1 vccd1 vccd1 _5208_/B sky130_fd_sc_hd__nand2_4
XFILLER_69_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5138_ _5138_/A _5138_/B vssd1 vssd1 vccd1 vccd1 _5138_/Y sky130_fd_sc_hd__nand2_2
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5069_ _5080_/B vssd1 vssd1 vccd1 vccd1 _5070_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4440_ _4267_/Y _4568_/A _3223_/B _5931_/A _4600_/A vssd1 vssd1 vccd1 vccd1 _4441_/C
+ sky130_fd_sc_hd__o2111ai_4
X_6110_ _6110_/A _6110_/B _6159_/A _6110_/D vssd1 vssd1 vccd1 vccd1 _6112_/B sky130_fd_sc_hd__nand4_1
X_4371_ _4182_/Y _4197_/Y _4368_/Y _4370_/Y vssd1 vssd1 vccd1 vccd1 _4371_/Y sky130_fd_sc_hd__o2bb2ai_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _3322_/A vssd1 vssd1 vccd1 vccd1 _4884_/A sky130_fd_sc_hd__clkbuf_2
X_6041_ _6041_/A _6041_/B vssd1 vssd1 vccd1 vccd1 _6041_/Y sky130_fd_sc_hd__nand2_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3897_/A vssd1 vssd1 vccd1 vccd1 _3414_/B sky130_fd_sc_hd__clkbuf_4
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _3184_/A _3229_/D _3310_/B _3184_/D vssd1 vssd1 vccd1 vccd1 _3242_/B sky130_fd_sc_hd__nand4_1
XFILLER_54_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5825_ _5852_/A _5825_/B _5852_/C _5825_/D vssd1 vssd1 vccd1 vccd1 _5825_/X sky130_fd_sc_hd__and4_1
XFILLER_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5756_ _5748_/X _5749_/Y _5751_/Y vssd1 vssd1 vccd1 vccd1 _5756_/Y sky130_fd_sc_hd__o21ai_1
X_5687_ _5590_/Y _5686_/Y _5609_/B vssd1 vssd1 vccd1 vccd1 _5744_/A sky130_fd_sc_hd__o21ai_1
X_4707_ _4703_/X _4704_/X _4705_/Y _4706_/Y vssd1 vssd1 vccd1 vccd1 _4988_/A sky130_fd_sc_hd__o211ai_4
X_4638_ _4641_/A _4469_/Y _4641_/B vssd1 vssd1 vccd1 vccd1 _4639_/C sky130_fd_sc_hd__o21ai_1
XFILLER_89_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4569_ _4569_/A vssd1 vssd1 vccd1 vccd1 _5065_/B sky130_fd_sc_hd__buf_4
XFILLER_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6239_ _6252_/A _6258_/A vssd1 vssd1 vccd1 vccd1 _6257_/A sky130_fd_sc_hd__nor2_1
XFILLER_49_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3940_ _4133_/B _3929_/Y _3985_/A _3985_/B vssd1 vssd1 vccd1 vccd1 _3973_/A sky130_fd_sc_hd__o211ai_2
XFILLER_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3871_ _5207_/A vssd1 vssd1 vccd1 vccd1 _4788_/A sky130_fd_sc_hd__buf_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5610_ _5590_/Y _5608_/X _5609_/Y vssd1 vssd1 vccd1 vccd1 _5611_/B sky130_fd_sc_hd__o21ai_4
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5541_ _5541_/A _5541_/B vssd1 vssd1 vccd1 vccd1 _5542_/B sky130_fd_sc_hd__nand2_1
X_5472_ _5303_/A _5303_/B _5297_/Y vssd1 vssd1 vccd1 vccd1 _5475_/B sky130_fd_sc_hd__o21a_1
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4423_ _4423_/A vssd1 vssd1 vccd1 vccd1 _5435_/A sky130_fd_sc_hd__clkbuf_4
X_4354_ input5/X vssd1 vssd1 vccd1 vccd1 _5299_/D sky130_fd_sc_hd__buf_2
XFILLER_86_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ _3293_/Y _3226_/A _3296_/Y vssd1 vssd1 vccd1 vccd1 _3305_/Y sky130_fd_sc_hd__o21ai_1
X_6024_ _6024_/A _6024_/B vssd1 vssd1 vccd1 vccd1 _6024_/Y sky130_fd_sc_hd__nand2_1
X_4285_ _4064_/X _4079_/Y _4071_/Y vssd1 vssd1 vccd1 vccd1 _4285_/Y sky130_fd_sc_hd__o21ai_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3236_ _3829_/B _5845_/A vssd1 vssd1 vccd1 vccd1 _3236_/Y sky130_fd_sc_hd__nand2_1
X_3167_ _3190_/A _3639_/A _3190_/C _3966_/B vssd1 vssd1 vccd1 vccd1 _3167_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_42_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5808_ _5808_/A _5808_/B vssd1 vssd1 vccd1 vccd1 _5808_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5739_ _5549_/C _5549_/A _5549_/B _5561_/C _5550_/A vssd1 vssd1 vccd1 vccd1 _5739_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4070_ _3891_/A _4064_/X _4067_/Y _4069_/Y vssd1 vssd1 vccd1 vccd1 _4070_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4972_ _4972_/A _4972_/B _4972_/C vssd1 vssd1 vccd1 vccd1 _4972_/Y sky130_fd_sc_hd__nand3_2
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3923_ _3902_/A _3902_/B _3918_/A vssd1 vssd1 vccd1 vccd1 _3923_/Y sky130_fd_sc_hd__a21oi_2
X_3854_ _3840_/X _3996_/B _3856_/A _3853_/Y _3849_/Y vssd1 vssd1 vccd1 vccd1 _4163_/B
+ sky130_fd_sc_hd__o221ai_4
X_3785_ _4708_/A _4238_/D vssd1 vssd1 vccd1 vccd1 _3787_/A sky130_fd_sc_hd__nand2_1
X_5524_ _5643_/A _5643_/B vssd1 vssd1 vccd1 vccd1 _5639_/A sky130_fd_sc_hd__nand2_1
X_5455_ _5288_/Y _5296_/D _5290_/Y vssd1 vssd1 vccd1 vccd1 _5457_/B sky130_fd_sc_hd__a21o_1
X_4406_ _4593_/A _4619_/B vssd1 vssd1 vccd1 vccd1 _4406_/Y sky130_fd_sc_hd__nand2_1
X_5386_ _5831_/B vssd1 vssd1 vccd1 vccd1 _5676_/A sky130_fd_sc_hd__buf_2
X_4337_ _4519_/A _4335_/A _4520_/A vssd1 vssd1 vccd1 vccd1 _4340_/B sky130_fd_sc_hd__a21o_1
XFILLER_59_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4268_ _4079_/Y _4267_/Y _4429_/A _4071_/B vssd1 vssd1 vccd1 vccd1 _4270_/A sky130_fd_sc_hd__o2bb2ai_1
X_6007_ _5927_/A _5927_/B _5927_/C vssd1 vssd1 vccd1 vccd1 _6007_/X sky130_fd_sc_hd__a21bo_1
X_3219_ _3256_/A vssd1 vssd1 vccd1 vccd1 _4025_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4199_ input5/X vssd1 vssd1 vccd1 vccd1 _4384_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3570_ _3472_/A _3472_/B _3477_/B _3477_/A vssd1 vssd1 vccd1 vccd1 _3570_/Y sky130_fd_sc_hd__a22oi_2
X_5240_ _5240_/A _5240_/B _5378_/B _5240_/D vssd1 vssd1 vccd1 vccd1 _5240_/X sky130_fd_sc_hd__and4_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5171_ _5175_/A _5175_/B _5171_/C _5171_/D vssd1 vssd1 vccd1 vccd1 _5172_/C sky130_fd_sc_hd__nand4_2
X_4122_ _4122_/A _4122_/B vssd1 vssd1 vccd1 vccd1 _4124_/B sky130_fd_sc_hd__nand2_2
X_4053_ _4054_/A _4054_/B _4054_/C vssd1 vssd1 vccd1 vccd1 _4053_/Y sky130_fd_sc_hd__a21oi_2
Xinput3 a[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4955_ _5132_/A _5532_/C _5532_/D _3783_/A vssd1 vssd1 vccd1 vccd1 _4955_/Y sky130_fd_sc_hd__a22oi_4
X_3906_ _3898_/X _3901_/X _3905_/X vssd1 vssd1 vccd1 vccd1 _4128_/A sky130_fd_sc_hd__o21ai_4
XFILLER_51_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4886_ _4885_/B _4885_/C _4885_/A vssd1 vssd1 vccd1 vccd1 _4886_/Y sky130_fd_sc_hd__a21oi_1
X_3837_ _3837_/A _3837_/B _3837_/C vssd1 vssd1 vccd1 vccd1 _3839_/B sky130_fd_sc_hd__nand3_2
X_3768_ _3414_/B _4936_/A _4238_/C _3418_/A vssd1 vssd1 vccd1 vccd1 _3768_/Y sky130_fd_sc_hd__a22oi_4
X_5507_ _5465_/C _4621_/C _5506_/X _6255_/A _5303_/B vssd1 vssd1 vccd1 vccd1 _5509_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_3_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3699_ _3699_/A _3699_/B vssd1 vssd1 vccd1 vccd1 _3699_/Y sky130_fd_sc_hd__nand2_1
X_5438_ _5464_/A _5465_/A vssd1 vssd1 vccd1 vccd1 _5438_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5369_ _5277_/Y _5367_/Y _5368_/Y vssd1 vssd1 vccd1 vccd1 _5483_/A sky130_fd_sc_hd__a21oi_1
XFILLER_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4740_ _4568_/B _4853_/A _3223_/B _5792_/B _4746_/A vssd1 vssd1 vccd1 vccd1 _4741_/C
+ sky130_fd_sc_hd__o2111ai_1
X_4671_ _4671_/A _4671_/B _4671_/C vssd1 vssd1 vccd1 vccd1 _4680_/D sky130_fd_sc_hd__nand3_2
X_3622_ _5037_/A vssd1 vssd1 vccd1 vccd1 _5401_/A sky130_fd_sc_hd__buf_4
X_3553_ _3280_/A _3474_/A _3419_/B _3676_/A _3552_/Y vssd1 vssd1 vccd1 vccd1 _3559_/A
+ sky130_fd_sc_hd__o221ai_4
X_6272_ _6247_/B _6247_/A _6267_/Y _6271_/Y vssd1 vssd1 vccd1 vccd1 _6273_/B sky130_fd_sc_hd__o211ai_2
X_3484_ _3484_/A _3484_/B vssd1 vssd1 vccd1 vccd1 _3584_/C sky130_fd_sc_hd__nand2_1
XFILLER_69_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5223_ _5223_/A vssd1 vssd1 vccd1 vccd1 _5808_/A sky130_fd_sc_hd__clkbuf_4
X_5154_ _5325_/A _5157_/B _5151_/Y _5153_/X vssd1 vssd1 vccd1 vccd1 _5159_/A sky130_fd_sc_hd__o2bb2ai_1
X_4105_ _4302_/A _4105_/B _5007_/A _5578_/A vssd1 vssd1 vccd1 vccd1 _4105_/Y sky130_fd_sc_hd__nand4_2
XFILLER_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5085_ _5085_/A _5104_/A vssd1 vssd1 vccd1 vccd1 _5278_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4036_ _3473_/Y _4372_/A _4025_/Y _4182_/A _4020_/Y vssd1 vssd1 vccd1 vccd1 _4036_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_71_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5987_ _5811_/A _6017_/A _5933_/C _6283_/C _5933_/A vssd1 vssd1 vccd1 vccd1 _5987_/Y
+ sky130_fd_sc_hd__o2111ai_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4938_ _4698_/Y _4929_/Y _4934_/Y _4937_/X vssd1 vssd1 vccd1 vccd1 _4938_/Y sky130_fd_sc_hd__a2bb2oi_4
X_4869_ _5087_/A _5087_/B _4868_/Y vssd1 vssd1 vccd1 vccd1 _4869_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5910_ _5914_/A _5914_/B _5914_/C _5914_/D vssd1 vssd1 vccd1 vccd1 _5911_/B sky130_fd_sc_hd__and4_1
XFILLER_19_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5841_ _3512_/X _6202_/B _5846_/B vssd1 vssd1 vccd1 vccd1 _5914_/B sky130_fd_sc_hd__o21ai_4
X_5772_ _5781_/A _5782_/A _5771_/X _5531_/Y vssd1 vssd1 vccd1 vccd1 _5773_/C sky130_fd_sc_hd__o2bb2ai_1
XFILLER_34_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4723_ _4721_/X _4722_/Y _4719_/Y _4712_/Y vssd1 vssd1 vccd1 vccd1 _4723_/X sky130_fd_sc_hd__o211a_2
X_4654_ _4647_/A _4498_/C _4648_/A vssd1 vssd1 vccd1 vccd1 _4661_/A sky130_fd_sc_hd__a21boi_4
X_3605_ _3607_/B _3607_/C _3607_/A vssd1 vssd1 vccd1 vccd1 _3605_/Y sky130_fd_sc_hd__a21oi_1
X_4585_ _4443_/Y _4575_/Y _4600_/B vssd1 vssd1 vccd1 vccd1 _4586_/C sky130_fd_sc_hd__o21ai_1
X_3536_ _3536_/A vssd1 vssd1 vccd1 vccd1 _4532_/A sky130_fd_sc_hd__clkbuf_2
X_6255_ _6255_/A _6255_/B _6255_/C _6283_/B vssd1 vssd1 vccd1 vccd1 _6260_/B sky130_fd_sc_hd__and4_1
XFILLER_88_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5206_ _5206_/A vssd1 vssd1 vccd1 vccd1 _5704_/A sky130_fd_sc_hd__buf_2
X_3467_ _3459_/Y _3462_/Y _3446_/X vssd1 vssd1 vccd1 vccd1 _3472_/A sky130_fd_sc_hd__o21ai_1
XFILLER_69_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6186_ _6222_/A _6187_/C _6187_/A vssd1 vssd1 vccd1 vccd1 _6190_/C sky130_fd_sc_hd__o21a_1
X_3398_ _3398_/A _3398_/B _3398_/C vssd1 vssd1 vccd1 vccd1 _3398_/X sky130_fd_sc_hd__and3_1
XFILLER_69_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5137_ _3350_/Y _4711_/C _5141_/B _5141_/C vssd1 vssd1 vccd1 vccd1 _5138_/B sky130_fd_sc_hd__o211ai_1
X_5068_ _5245_/A _5068_/B _5397_/B _5068_/D vssd1 vssd1 vccd1 vccd1 _5080_/B sky130_fd_sc_hd__nand4_4
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4019_ _4019_/A _5286_/A vssd1 vssd1 vccd1 vccd1 _4020_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4370_ _4182_/B _4529_/A _4366_/Y vssd1 vssd1 vccd1 vccd1 _4370_/Y sky130_fd_sc_hd__o21ai_1
X_3321_ _5663_/A vssd1 vssd1 vccd1 vccd1 _5905_/A sky130_fd_sc_hd__buf_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6040_/A _6101_/A _6041_/B vssd1 vssd1 vccd1 vccd1 _6047_/A sky130_fd_sc_hd__nand3_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3551_/A vssd1 vssd1 vccd1 vccd1 _3677_/A sky130_fd_sc_hd__clkbuf_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _3829_/B _3229_/D _3184_/D _3184_/A vssd1 vssd1 vccd1 vccd1 _3242_/A sky130_fd_sc_hd__a22o_1
XFILLER_78_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5824_ _6077_/B vssd1 vssd1 vccd1 vccd1 _5825_/D sky130_fd_sc_hd__buf_2
X_5755_ _5693_/X _5746_/Y _5753_/Y _5754_/X vssd1 vssd1 vccd1 vccd1 _5884_/A sky130_fd_sc_hd__o211ai_4
X_5686_ _5686_/A _5686_/B vssd1 vssd1 vccd1 vccd1 _5686_/Y sky130_fd_sc_hd__nand2_1
X_4706_ _4703_/X _4698_/Y _4700_/Y vssd1 vssd1 vccd1 vccd1 _4706_/Y sky130_fd_sc_hd__o21ai_2
X_4637_ _4634_/Y _4635_/X _4643_/A _4643_/B vssd1 vssd1 vccd1 vccd1 _4639_/B sky130_fd_sc_hd__o211ai_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4568_ _4568_/A _4568_/B vssd1 vssd1 vccd1 vccd1 _4576_/B sky130_fd_sc_hd__nand2_2
X_3519_ _5833_/B vssd1 vssd1 vccd1 vccd1 _5994_/A sky130_fd_sc_hd__clkbuf_4
X_4499_ _4499_/A _4499_/B _4499_/C vssd1 vssd1 vccd1 vccd1 _4502_/B sky130_fd_sc_hd__nand3_1
X_6238_ _6236_/X _6208_/A _6234_/X _6235_/Y vssd1 vssd1 vccd1 vccd1 _6258_/A sky130_fd_sc_hd__a211oi_4
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6169_ _6170_/B _6072_/C _6170_/D _6203_/A vssd1 vssd1 vccd1 vccd1 _6171_/B sky130_fd_sc_hd__a22oi_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3870_ _3870_/A vssd1 vssd1 vccd1 vccd1 _4700_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5540_ _5697_/A vssd1 vssd1 vccd1 vccd1 _5540_/X sky130_fd_sc_hd__buf_2
X_5471_ _5471_/A _5471_/B _5471_/C vssd1 vssd1 vccd1 vccd1 _5634_/A sky130_fd_sc_hd__nand3_4
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4422_ _4422_/A _4422_/B _4422_/C vssd1 vssd1 vccd1 vccd1 _4422_/X sky130_fd_sc_hd__and3_1
X_4353_ _4193_/A _5532_/C _5532_/D _3960_/B vssd1 vssd1 vccd1 vccd1 _4680_/A sky130_fd_sc_hd__a22o_2
X_4284_ _4284_/A _4284_/B _4284_/C vssd1 vssd1 vccd1 vccd1 _4284_/X sky130_fd_sc_hd__and3_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3304_ _3345_/B _3287_/X _3345_/A vssd1 vssd1 vccd1 vccd1 _3304_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6023_ _6091_/A _6023_/B _6023_/C vssd1 vssd1 vccd1 vccd1 _6024_/B sky130_fd_sc_hd__nand3_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _5678_/A vssd1 vssd1 vccd1 vccd1 _5845_/A sky130_fd_sc_hd__buf_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3166_ _3803_/A vssd1 vssd1 vccd1 vccd1 _3639_/A sky130_fd_sc_hd__buf_2
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5807_ _5811_/B _6077_/A _5809_/A _5712_/A _4829_/A vssd1 vssd1 vccd1 vccd1 _5807_/Y
+ sky130_fd_sc_hd__a32oi_4
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3999_ _3999_/A _3999_/B vssd1 vssd1 vccd1 vccd1 _4161_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5738_ _5735_/Y _5736_/Y _5737_/Y vssd1 vssd1 vccd1 vccd1 _5738_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5669_ _5669_/A _5842_/A vssd1 vssd1 vccd1 vccd1 _5832_/A sky130_fd_sc_hd__nand2_1
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4971_ _5175_/A _4988_/D _4971_/C vssd1 vssd1 vccd1 vccd1 _4984_/B sky130_fd_sc_hd__and3_1
XFILLER_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3922_ _3780_/X _3764_/A _3757_/X _3752_/X vssd1 vssd1 vccd1 vccd1 _3928_/A sky130_fd_sc_hd__o2bb2ai_1
X_3853_ _3853_/A _3856_/B vssd1 vssd1 vccd1 vccd1 _3853_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3784_ _3676_/A _3676_/B _3783_/Y vssd1 vssd1 vccd1 vccd1 _3784_/Y sky130_fd_sc_hd__a21oi_1
X_5523_ _5523_/A _5523_/B vssd1 vssd1 vccd1 vccd1 _5523_/X sky130_fd_sc_hd__xor2_4
X_5454_ _5454_/A _5454_/B vssd1 vssd1 vccd1 vccd1 _5457_/A sky130_fd_sc_hd__nand2_1
X_4405_ _3620_/C _5532_/A _4236_/B _5399_/A vssd1 vssd1 vccd1 vccd1 _4405_/Y sky130_fd_sc_hd__a22oi_2
X_5385_ _5681_/A vssd1 vssd1 vccd1 vccd1 _6236_/B sky130_fd_sc_hd__inv_2
X_4336_ _4520_/A _4519_/A _4519_/B vssd1 vssd1 vccd1 vccd1 _4340_/A sky130_fd_sc_hd__nand3_1
XFILLER_86_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4267_ _4855_/A _5207_/B vssd1 vssd1 vccd1 vccd1 _4267_/Y sky130_fd_sc_hd__nand2_2
X_6006_ _6006_/A _6134_/C _6132_/C _6006_/D vssd1 vssd1 vccd1 vccd1 _6006_/X sky130_fd_sc_hd__and4_1
X_3218_ _3218_/A _3458_/B _3555_/A _3783_/A vssd1 vssd1 vccd1 vccd1 _3229_/B sky130_fd_sc_hd__nand4_2
X_4198_ _4186_/Y _4189_/Y _4196_/Y _4197_/Y _4023_/Y vssd1 vssd1 vccd1 vccd1 _4198_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3149_ _3310_/B vssd1 vssd1 vccd1 vccd1 _4832_/C sky130_fd_sc_hd__buf_2
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5170_ _5176_/A _5170_/B vssd1 vssd1 vccd1 vccd1 _5172_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4121_ _4220_/A _4135_/B _4127_/C vssd1 vssd1 vccd1 vccd1 _4122_/B sky130_fd_sc_hd__nand3_1
XFILLER_68_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4052_ _4052_/A vssd1 vssd1 vccd1 vccd1 _4054_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 a[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
XFILLER_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4954_ _4698_/Y _4929_/Y _4952_/X _4953_/Y vssd1 vssd1 vccd1 vccd1 _4954_/Y sky130_fd_sc_hd__o211ai_4
X_3905_ _4880_/A _3543_/B _3918_/B _3918_/C vssd1 vssd1 vccd1 vccd1 _3905_/X sky130_fd_sc_hd__a22o_1
XFILLER_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4885_ _4885_/A _4885_/B _4885_/C vssd1 vssd1 vccd1 vccd1 _4885_/X sky130_fd_sc_hd__and3_1
X_3836_ _3836_/A _3836_/B vssd1 vssd1 vccd1 vccd1 _3847_/B sky130_fd_sc_hd__nand2_1
X_3767_ _4693_/A vssd1 vssd1 vccd1 vccd1 _4238_/C sky130_fd_sc_hd__buf_4
X_5506_ _5506_/A vssd1 vssd1 vccd1 vccd1 _5506_/X sky130_fd_sc_hd__clkbuf_4
X_3698_ _3558_/A _3560_/B _3558_/B vssd1 vssd1 vccd1 vccd1 _3719_/A sky130_fd_sc_hd__a21boi_1
X_5437_ _5437_/A _5437_/B vssd1 vssd1 vccd1 vccd1 _5465_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5368_ _5277_/B _5277_/C _5277_/A vssd1 vssd1 vccd1 vccd1 _5368_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4319_ _4322_/A _4322_/B _4224_/X _4318_/Y vssd1 vssd1 vccd1 vccd1 _4323_/B sky130_fd_sc_hd__o2bb2ai_1
X_5299_ _5299_/A _5299_/B _5299_/C _5299_/D vssd1 vssd1 vccd1 vccd1 _5514_/A sky130_fd_sc_hd__nand4_4
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4670_ _4663_/A _4663_/B _4669_/Y vssd1 vssd1 vccd1 vccd1 _4671_/C sky130_fd_sc_hd__a21o_1
X_3621_ _3473_/Y _3512_/X _3806_/A _3630_/B vssd1 vssd1 vccd1 vccd1 _3625_/B sky130_fd_sc_hd__o211ai_2
X_3552_ _3552_/A _3611_/A vssd1 vssd1 vccd1 vccd1 _3552_/Y sky130_fd_sc_hd__nand2_1
X_6271_ _6271_/A _6271_/B vssd1 vssd1 vccd1 vccd1 _6271_/Y sky130_fd_sc_hd__nand2_1
X_3483_ _3483_/A _3483_/B vssd1 vssd1 vccd1 vccd1 _3484_/B sky130_fd_sc_hd__nand2_1
X_5222_ _5222_/A vssd1 vssd1 vccd1 vccd1 _5281_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5153_ _4965_/X _5152_/X _5163_/B _5145_/A vssd1 vssd1 vccd1 vccd1 _5153_/X sky130_fd_sc_hd__o211a_1
X_4104_ _4700_/A _4945_/A _4788_/A _4238_/D vssd1 vssd1 vccd1 vccd1 _4105_/B sky130_fd_sc_hd__nand4_4
X_5084_ _5084_/A _5084_/B _5084_/C vssd1 vssd1 vccd1 vccd1 _5104_/A sky130_fd_sc_hd__nand3_1
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4035_ input3/X vssd1 vssd1 vccd1 vccd1 _4372_/A sky130_fd_sc_hd__clkinv_2
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5986_ _6079_/A _5986_/B vssd1 vssd1 vccd1 vccd1 _6017_/A sky130_fd_sc_hd__nand2_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4937_ _4933_/X _4935_/Y _4936_/Y vssd1 vssd1 vccd1 vccd1 _4937_/X sky130_fd_sc_hd__a21o_1
XANTENNA_20 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4868_ _4868_/A _5068_/D vssd1 vssd1 vccd1 vccd1 _4868_/Y sky130_fd_sc_hd__nand2_1
X_3819_ _3819_/A _3819_/B _3819_/C vssd1 vssd1 vccd1 vccd1 _3822_/C sky130_fd_sc_hd__nand3_4
X_4799_ _4607_/B _4794_/Y _4795_/Y vssd1 vssd1 vccd1 vccd1 _4803_/A sky130_fd_sc_hd__o21ai_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5840_ _5840_/A _5840_/B _5840_/C vssd1 vssd1 vccd1 vccd1 _5840_/Y sky130_fd_sc_hd__nand3_2
X_5771_ _3669_/X _4674_/X _5437_/B _5534_/Y vssd1 vssd1 vccd1 vccd1 _5771_/X sky130_fd_sc_hd__o22a_1
XFILLER_61_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4722_ _4722_/A _4722_/B vssd1 vssd1 vccd1 vccd1 _4722_/Y sky130_fd_sc_hd__nand2_1
X_4653_ _4653_/A vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__clkbuf_4
X_3604_ _3366_/Y _3369_/Y _3362_/Y _3410_/A vssd1 vssd1 vccd1 vccd1 _3607_/A sky130_fd_sc_hd__a211o_2
X_4584_ _4581_/A _4731_/A _5240_/B _5701_/B _4576_/B vssd1 vssd1 vccd1 vccd1 _4586_/B
+ sky130_fd_sc_hd__o2111ai_1
X_3535_ _3441_/X _4417_/A _3564_/A _3564_/B vssd1 vssd1 vccd1 vccd1 _3535_/Y sky130_fd_sc_hd__o211ai_1
X_6254_ _6255_/B _6255_/C _6283_/B _5967_/X vssd1 vssd1 vccd1 vccd1 _6260_/A sky130_fd_sc_hd__a22oi_2
X_3466_ _3459_/Y _3462_/Y _3446_/X _3465_/Y vssd1 vssd1 vccd1 vccd1 _3478_/A sky130_fd_sc_hd__o211ai_2
X_5205_ _4236_/A _5701_/B _4875_/B _5250_/A vssd1 vssd1 vccd1 vccd1 _5205_/X sky130_fd_sc_hd__o2bb2a_1
X_6185_ _5506_/X _5967_/X _5825_/D _6072_/C _6138_/B vssd1 vssd1 vccd1 vccd1 _6187_/A
+ sky130_fd_sc_hd__a41oi_4
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3397_ _3598_/A _3315_/C _3598_/C _3396_/X vssd1 vssd1 vccd1 vccd1 _3397_/X sky130_fd_sc_hd__o31a_1
X_5136_ _5136_/A vssd1 vssd1 vccd1 vccd1 _5141_/C sky130_fd_sc_hd__buf_2
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5067_ _5067_/A _5067_/B vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4018_ _4025_/A _5539_/A vssd1 vssd1 vccd1 vccd1 _4020_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5969_ _6058_/A _5969_/B _5969_/C vssd1 vssd1 vccd1 vccd1 _5971_/A sky130_fd_sc_hd__nand3_1
XFILLER_75_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3320_ _5209_/A vssd1 vssd1 vccd1 vccd1 _5663_/A sky130_fd_sc_hd__buf_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3772_/A vssd1 vssd1 vccd1 vccd1 _3551_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3182_ _3639_/A _3179_/C _5006_/A _3218_/A vssd1 vssd1 vccd1 vccd1 _3184_/A sky130_fd_sc_hd__a22o_1
XFILLER_78_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5823_ _5823_/A vssd1 vssd1 vccd1 vccd1 _5944_/B sky130_fd_sc_hd__inv_2
XFILLER_22_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5754_ _5625_/A _5625_/B _5625_/D _5619_/Y vssd1 vssd1 vccd1 vccd1 _5754_/X sky130_fd_sc_hd__a31o_1
X_5685_ _5673_/Y _5675_/X _5684_/Y vssd1 vssd1 vccd1 vccd1 _5685_/X sky130_fd_sc_hd__a21bo_1
X_4705_ _4690_/Y _4691_/Y _4530_/Y vssd1 vssd1 vccd1 vccd1 _4705_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4636_ _4636_/A vssd1 vssd1 vccd1 vccd1 _4643_/B sky130_fd_sc_hd__buf_2
XFILLER_1_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4567_ _5045_/A _4863_/A vssd1 vssd1 vccd1 vccd1 _4568_/B sky130_fd_sc_hd__nand2_1
X_3518_ _5404_/B vssd1 vssd1 vccd1 vccd1 _5833_/B sky130_fd_sc_hd__buf_2
X_4498_ _4647_/A _4648_/A _4498_/C vssd1 vssd1 vccd1 vccd1 _4499_/C sky130_fd_sc_hd__nand3_1
X_6237_ _6234_/X _6235_/Y _6236_/X _6208_/A vssd1 vssd1 vccd1 vccd1 _6252_/A sky130_fd_sc_hd__o211a_1
X_3449_ _5603_/A _3448_/X _3439_/A vssd1 vssd1 vccd1 vccd1 _3452_/B sky130_fd_sc_hd__o21ai_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6132_/B _6132_/Y _6165_/X _6166_/Y vssd1 vssd1 vccd1 vccd1 _6199_/A sky130_fd_sc_hd__a211o_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5119_ _5119_/A _5123_/A _5286_/A _5119_/D vssd1 vssd1 vccd1 vccd1 _5128_/B sky130_fd_sc_hd__nand4_4
XFILLER_84_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6099_ _6101_/A _6151_/A _6100_/B vssd1 vssd1 vccd1 vccd1 _6104_/B sky130_fd_sc_hd__nand3b_1
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5470_ _5026_/Y _5281_/B _5469_/X _5432_/Y vssd1 vssd1 vccd1 vccd1 _5471_/C sky130_fd_sc_hd__a31oi_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4421_ _4232_/Y _4230_/Y _4238_/Y _4414_/X _4420_/X vssd1 vssd1 vccd1 vccd1 _4489_/A
+ sky130_fd_sc_hd__o2111ai_4
X_4352_ input5/X vssd1 vssd1 vccd1 vccd1 _5532_/D sky130_fd_sc_hd__clkbuf_4
X_4283_ _4298_/C _4298_/D vssd1 vssd1 vccd1 vccd1 _4283_/Y sky130_fd_sc_hd__nand2_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3303_ _3240_/A _3240_/C _3240_/B vssd1 vssd1 vccd1 vccd1 _3309_/A sky130_fd_sc_hd__a21boi_1
X_6022_ _6091_/A _6091_/B _6023_/C vssd1 vssd1 vccd1 vccd1 _6022_/Y sky130_fd_sc_hd__a21oi_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _4235_/B vssd1 vssd1 vccd1 vccd1 _5678_/A sky130_fd_sc_hd__buf_2
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3165_ _3190_/A _4827_/A _3190_/C _3310_/B vssd1 vssd1 vccd1 vccd1 _3165_/X sky130_fd_sc_hd__and4_1
XFILLER_27_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5806_ _6020_/C _6170_/A _5811_/B vssd1 vssd1 vccd1 vccd1 _5806_/X sky130_fd_sc_hd__a21o_1
X_3998_ _3998_/A _4166_/A _3998_/C _3998_/D vssd1 vssd1 vccd1 vccd1 _4004_/A sky130_fd_sc_hd__or4_1
X_5737_ _5729_/A _5729_/B _5728_/A _5728_/B vssd1 vssd1 vccd1 vccd1 _5737_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_22_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5668_ _5604_/A _5592_/Y _5604_/B vssd1 vssd1 vccd1 vccd1 _5826_/B sky130_fd_sc_hd__o21ai_1
X_4619_ _4788_/A _4619_/B _5575_/A _5037_/B vssd1 vssd1 vccd1 vccd1 _4621_/B sky130_fd_sc_hd__nand4_4
X_5599_ _5599_/A vssd1 vssd1 vccd1 vccd1 _6235_/B sky130_fd_sc_hd__buf_2
XFILLER_89_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _5175_/A _4988_/D _4971_/C vssd1 vssd1 vccd1 vccd1 _4984_/A sky130_fd_sc_hd__a21oi_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3921_ _3938_/A _3938_/B _3936_/A vssd1 vssd1 vccd1 vccd1 _4133_/B sky130_fd_sc_hd__o21ai_2
X_3852_ _3998_/C _3852_/B vssd1 vssd1 vccd1 vccd1 _4163_/A sky130_fd_sc_hd__nand2_1
X_5522_ _5980_/A _5980_/B _5521_/Y vssd1 vssd1 vccd1 vccd1 _5523_/B sky130_fd_sc_hd__a21oi_4
X_3783_ _3783_/A _5248_/A vssd1 vssd1 vccd1 vccd1 _3783_/Y sky130_fd_sc_hd__nand2_1
X_5453_ _5453_/A _5453_/B vssd1 vssd1 vccd1 vccd1 _5454_/B sky130_fd_sc_hd__nor2_1
X_5384_ _5677_/A vssd1 vssd1 vccd1 vccd1 _5681_/A sky130_fd_sc_hd__clkbuf_2
X_4404_ _4931_/A vssd1 vssd1 vccd1 vccd1 _5532_/A sky130_fd_sc_hd__buf_2
X_4335_ _4335_/A vssd1 vssd1 vccd1 vccd1 _4519_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4266_ _3894_/A _4261_/Y _4057_/X _4429_/A _4277_/A vssd1 vssd1 vccd1 vccd1 _4266_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_86_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6005_ _6205_/C _5825_/D _6006_/D _6006_/A vssd1 vssd1 vccd1 vccd1 _6005_/Y sky130_fd_sc_hd__a22oi_2
X_3217_ _3866_/A vssd1 vssd1 vccd1 vccd1 _3783_/A sky130_fd_sc_hd__clkbuf_4
X_4197_ _4197_/A _4197_/B vssd1 vssd1 vccd1 vccd1 _4197_/Y sky130_fd_sc_hd__nand2_2
X_3148_ _3966_/B vssd1 vssd1 vccd1 vccd1 _3310_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4120_ _4211_/A vssd1 vssd1 vccd1 vccd1 _4135_/B sky130_fd_sc_hd__clkbuf_2
X_4051_ _4051_/A vssd1 vssd1 vccd1 vccd1 _4054_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput5 a[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4953_ _4928_/X _5124_/A _5347_/A _4179_/X _4933_/X vssd1 vssd1 vccd1 vccd1 _4953_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_3904_ _5245_/A _5068_/B _5119_/A _4693_/A vssd1 vssd1 vccd1 vccd1 _3918_/C sky130_fd_sc_hd__nand4_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4884_ _4884_/A _4884_/B vssd1 vssd1 vccd1 vccd1 _4885_/A sky130_fd_sc_hd__nand2_2
X_3835_ _3835_/A _3835_/B vssd1 vssd1 vccd1 vccd1 _3836_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3766_ _3766_/A vssd1 vssd1 vccd1 vccd1 _4693_/A sky130_fd_sc_hd__buf_2
X_5505_ _5509_/C vssd1 vssd1 vccd1 vccd1 _5643_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5436_ _5436_/A _5436_/B vssd1 vssd1 vccd1 vccd1 _5437_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3697_ _3639_/X _3641_/X _3691_/X _3625_/Y vssd1 vssd1 vccd1 vccd1 _3697_/X sky130_fd_sc_hd__o211a_1
X_5367_ _5367_/A _5367_/B vssd1 vssd1 vccd1 vccd1 _5367_/Y sky130_fd_sc_hd__nand2_1
X_5298_ _5289_/Y _5293_/Y _5297_/Y vssd1 vssd1 vccd1 vccd1 _5304_/A sky130_fd_sc_hd__o21ai_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4318_ _4313_/B _4313_/C _4224_/C vssd1 vssd1 vccd1 vccd1 _4318_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4249_ _4302_/C _4302_/D _4250_/C vssd1 vssd1 vccd1 vccd1 _4249_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3620_ _4355_/A _4540_/B _3620_/C _5399_/A vssd1 vssd1 vccd1 vccd1 _3630_/B sky130_fd_sc_hd__nand4_2
X_3551_ _3551_/A _3867_/A vssd1 vssd1 vccd1 vccd1 _3611_/A sky130_fd_sc_hd__nand2_1
X_6270_ _6275_/C vssd1 vssd1 vccd1 vccd1 _6271_/B sky130_fd_sc_hd__inv_2
X_3482_ _3482_/A vssd1 vssd1 vccd1 vccd1 _3593_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5221_ _5222_/A _5271_/A _5219_/X _5220_/Y vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__o2bb2a_1
X_5152_ _4957_/X _4955_/Y _4959_/Y _4954_/Y vssd1 vssd1 vccd1 vccd1 _5152_/X sky130_fd_sc_hd__o211a_1
X_4103_ _4103_/A _4103_/B vssd1 vssd1 vccd1 vccd1 _4302_/A sky130_fd_sc_hd__nand2_2
X_5083_ _5078_/Y _5080_/X _5081_/X _5082_/Y _5095_/B vssd1 vssd1 vccd1 vccd1 _5084_/C
+ sky130_fd_sc_hd__o221ai_1
XFILLER_37_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4034_ _4177_/A _4177_/B _4177_/C vssd1 vssd1 vccd1 vccd1 _4048_/B sky130_fd_sc_hd__nand3_4
XFILLER_24_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5985_ _5983_/Y _5982_/B _5984_/X vssd1 vssd1 vccd1 vccd1 _6060_/A sky130_fd_sc_hd__a21bo_1
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4936_ _4936_/A _4936_/B vssd1 vssd1 vccd1 vccd1 _4936_/Y sky130_fd_sc_hd__nand2_2
XANTENNA_10 _5897_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _5982_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4867_ _3894_/A _5376_/A _4860_/X _5046_/A _5087_/A vssd1 vssd1 vccd1 vccd1 _4867_/Y
+ sky130_fd_sc_hd__o221ai_1
X_3818_ _3687_/A _3690_/Y _3720_/C vssd1 vssd1 vccd1 vccd1 _3837_/B sky130_fd_sc_hd__o21ai_4
XFILLER_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4798_ _4607_/B _4794_/Y _4795_/Y _4797_/Y vssd1 vssd1 vccd1 vccd1 _4798_/Y sky130_fd_sc_hd__o211ai_4
X_3749_ _4852_/A _4738_/A _4068_/A _4065_/A vssd1 vssd1 vccd1 vccd1 _3755_/B sky130_fd_sc_hd__nand4_4
X_5419_ _5420_/A _5254_/B _5256_/A vssd1 vssd1 vccd1 vccd1 _5419_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_87_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5770_ _5781_/A _5782_/A _5781_/B vssd1 vssd1 vccd1 vccd1 _5773_/B sky130_fd_sc_hd__nand3_1
XFILLER_61_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4721_ _4703_/X _4704_/X _4705_/Y _4706_/Y vssd1 vssd1 vccd1 vccd1 _4721_/X sky130_fd_sc_hd__o211a_2
X_4652_ _4652_/A _4652_/B _4652_/C vssd1 vssd1 vccd1 vccd1 _4653_/A sky130_fd_sc_hd__nand3_2
Xinput30 b[5] vssd1 vssd1 vccd1 vccd1 _3437_/A sky130_fd_sc_hd__clkbuf_2
X_3603_ _3586_/A _3586_/B _3586_/C _3857_/B _3857_/C vssd1 vssd1 vccd1 vccd1 _3603_/Y
+ sky130_fd_sc_hd__a32oi_4
X_4583_ _4873_/B vssd1 vssd1 vccd1 vccd1 _5701_/B sky130_fd_sc_hd__buf_2
X_3534_ _3657_/B vssd1 vssd1 vccd1 vccd1 _3564_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6253_ _6253_/A vssd1 vssd1 vccd1 vccd1 _6283_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3465_ _3465_/A _3465_/B vssd1 vssd1 vccd1 vccd1 _3465_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5204_ _3414_/B _5065_/B _5575_/B _3418_/A vssd1 vssd1 vccd1 vccd1 _5204_/Y sky130_fd_sc_hd__a22oi_4
X_6184_ _6183_/A _6183_/B _6182_/X vssd1 vssd1 vccd1 vccd1 _6187_/C sky130_fd_sc_hd__o21ba_1
X_3396_ _3598_/A _3315_/C _3597_/A _3395_/X vssd1 vssd1 vccd1 vccd1 _3396_/X sky130_fd_sc_hd__a2bb2o_1
X_5135_ _5141_/B _5136_/A _5141_/A vssd1 vssd1 vccd1 vccd1 _5138_/A sky130_fd_sc_hd__a21o_1
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5066_ _5066_/A _5570_/A vssd1 vssd1 vccd1 vccd1 _5067_/B sky130_fd_sc_hd__nand2_1
X_4017_ input2/X vssd1 vssd1 vccd1 vccd1 _5539_/A sky130_fd_sc_hd__buf_2
XFILLER_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5968_ _5933_/C _6020_/C _5506_/X _5967_/X _5812_/X vssd1 vssd1 vccd1 vccd1 _5969_/C
+ sky130_fd_sc_hd__a41o_1
X_4919_ _4922_/A _5100_/A _5100_/B vssd1 vssd1 vccd1 vccd1 _4919_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5899_ _5881_/X _5898_/Y _5872_/Y vssd1 vssd1 vccd1 vccd1 _5966_/C sky130_fd_sc_hd__o21ai_1
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3473_/A vssd1 vssd1 vccd1 vccd1 _3960_/B sky130_fd_sc_hd__clkbuf_4
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _3555_/A vssd1 vssd1 vccd1 vccd1 _5006_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5822_ _5944_/A _5945_/A vssd1 vssd1 vccd1 vccd1 _5822_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5753_ _5693_/X _5747_/Y _5752_/X vssd1 vssd1 vccd1 vccd1 _5753_/Y sky130_fd_sc_hd__o21ai_1
X_4704_ _3714_/D _4625_/A _5919_/A _6009_/A _4700_/Y vssd1 vssd1 vccd1 vccd1 _4704_/X
+ sky130_fd_sc_hd__a41o_1
X_5684_ _5840_/B _5684_/B vssd1 vssd1 vccd1 vccd1 _5684_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4635_ _4635_/A _4635_/B _4635_/C vssd1 vssd1 vccd1 vccd1 _4635_/X sky130_fd_sc_hd__and3_1
X_4566_ _4578_/A vssd1 vssd1 vccd1 vccd1 _4863_/A sky130_fd_sc_hd__clkbuf_2
X_3517_ _3730_/A _3522_/A _3402_/Y _3498_/A vssd1 vssd1 vccd1 vccd1 _3576_/A sky130_fd_sc_hd__o2bb2ai_2
XFILLER_1_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4497_ _4322_/A _4321_/A _4321_/B _4348_/Y vssd1 vssd1 vccd1 vccd1 _4499_/B sky130_fd_sc_hd__a31oi_1
X_6236_ _6236_/A _6236_/B _6236_/C vssd1 vssd1 vccd1 vccd1 _6236_/X sky130_fd_sc_hd__or3_1
X_3448_ _3448_/A vssd1 vssd1 vccd1 vccd1 _3448_/X sky130_fd_sc_hd__clkbuf_4
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6165_/X _6166_/Y _6132_/B _6132_/Y vssd1 vssd1 vccd1 vccd1 _6173_/A sky130_fd_sc_hd__o211ai_2
X_3379_ _3376_/Y _3360_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3381_/B sky130_fd_sc_hd__a21o_1
XFILLER_94_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _5299_/B _5288_/B vssd1 vssd1 vccd1 vccd1 _5120_/A sky130_fd_sc_hd__nand2_1
X_6098_ _6097_/A _6149_/B _6097_/C vssd1 vssd1 vccd1 vccd1 _6100_/B sky130_fd_sc_hd__a21o_1
XFILLER_57_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5049_ _5245_/B vssd1 vssd1 vccd1 vccd1 _5599_/A sky130_fd_sc_hd__inv_2
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4420_ _4420_/A vssd1 vssd1 vccd1 vccd1 _4420_/X sky130_fd_sc_hd__clkbuf_2
X_4351_ input4/X vssd1 vssd1 vccd1 vccd1 _5532_/C sky130_fd_sc_hd__buf_2
X_4282_ _4298_/A _4298_/B vssd1 vssd1 vccd1 vccd1 _4294_/C sky130_fd_sc_hd__nand2_2
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3302_ _3302_/A _3302_/B _3302_/C vssd1 vssd1 vccd1 vccd1 _3312_/A sky130_fd_sc_hd__nand3_1
X_6021_ _6021_/A _6110_/B vssd1 vssd1 vccd1 vccd1 _6023_/C sky130_fd_sc_hd__or2b_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _5065_/A vssd1 vssd1 vccd1 vccd1 _4235_/B sky130_fd_sc_hd__clkbuf_4
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3164_ _3791_/C vssd1 vssd1 vccd1 vccd1 _4827_/A sky130_fd_sc_hd__buf_2
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5805_ _5805_/A _5805_/B vssd1 vssd1 vccd1 vccd1 _5811_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3997_ _4163_/C vssd1 vssd1 vccd1 vccd1 _3998_/D sky130_fd_sc_hd__inv_2
X_5736_ _5588_/A _5588_/B _5588_/C _5608_/A vssd1 vssd1 vccd1 vccd1 _5736_/Y sky130_fd_sc_hd__a31oi_1
X_5667_ _4422_/B _6010_/B _5852_/A _5825_/B vssd1 vssd1 vccd1 vccd1 _5826_/A sky130_fd_sc_hd__a22o_1
X_4618_ _4618_/A _4618_/B vssd1 vssd1 vccd1 vccd1 _4621_/A sky130_fd_sc_hd__nand2_4
X_5598_ _5598_/A _5598_/B vssd1 vssd1 vccd1 vccd1 _5661_/A sky130_fd_sc_hd__nand2_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4549_ _4366_/Y _4368_/Y _4531_/Y _4548_/X _4363_/Y vssd1 vssd1 vccd1 vccd1 _4549_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6219_ _6219_/A _6219_/B _6219_/C vssd1 vssd1 vccd1 vccd1 _6220_/B sky130_fd_sc_hd__and3_1
XFILLER_89_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3920_ _3920_/A _3920_/B _3920_/C vssd1 vssd1 vccd1 vccd1 _3936_/A sky130_fd_sc_hd__nand3_2
XFILLER_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3851_ _3853_/A _3998_/A _3856_/B vssd1 vssd1 vccd1 vccd1 _3852_/B sky130_fd_sc_hd__a21o_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3782_ _3819_/A _3819_/B _3819_/C vssd1 vssd1 vccd1 vccd1 _3782_/X sky130_fd_sc_hd__and3_1
X_5521_ _5519_/X _5520_/X _5518_/C _5192_/Y vssd1 vssd1 vccd1 vccd1 _5521_/Y sky130_fd_sc_hd__o22ai_4
X_5452_ _5291_/X _5542_/A _5445_/Y vssd1 vssd1 vccd1 vccd1 _5454_/A sky130_fd_sc_hd__o21ai_1
X_4403_ _4411_/A _4411_/B _4402_/Y vssd1 vssd1 vccd1 vccd1 _4630_/B sky130_fd_sc_hd__o21ai_2
X_5383_ _5383_/A _5383_/B _5383_/C vssd1 vssd1 vccd1 vccd1 _5612_/A sky130_fd_sc_hd__nand3_4
X_4334_ _4334_/A _4334_/B _4334_/C vssd1 vssd1 vccd1 vccd1 _4335_/A sky130_fd_sc_hd__nand3_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6004_ _6004_/A _6004_/B vssd1 vssd1 vccd1 vccd1 _6006_/A sky130_fd_sc_hd__nand2_1
X_4265_ _4855_/B _5029_/B _4873_/B _4855_/A vssd1 vssd1 vccd1 vccd1 _4277_/A sky130_fd_sc_hd__a22o_1
XFILLER_67_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3216_ _3356_/A vssd1 vssd1 vccd1 vccd1 _3866_/A sky130_fd_sc_hd__clkbuf_2
X_4196_ _4363_/A _5794_/A _6009_/A _3555_/A vssd1 vssd1 vccd1 vccd1 _4196_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3147_ _4186_/A vssd1 vssd1 vccd1 vccd1 _3966_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_94_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5719_ _5719_/A _6137_/B _5719_/C _5719_/D vssd1 vssd1 vccd1 vccd1 _5733_/B sky130_fd_sc_hd__nand4_1
XFILLER_6_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4050_ _3981_/Y _4045_/Y _4048_/Y _4049_/X vssd1 vssd1 vccd1 vccd1 _4051_/A sky130_fd_sc_hd__o211ai_4
Xinput6 a[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_2
XFILLER_64_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4952_ _5347_/A _4038_/B _4933_/X _4935_/Y vssd1 vssd1 vccd1 vccd1 _4952_/X sky130_fd_sc_hd__a22o_1
X_3903_ _3903_/A vssd1 vssd1 vccd1 vccd1 _5119_/A sky130_fd_sc_hd__clkbuf_4
X_4883_ _4865_/Y _4871_/X _4879_/Y _4882_/X vssd1 vssd1 vccd1 vccd1 _4893_/A sky130_fd_sc_hd__o2bb2ai_1
X_3834_ _3821_/X _3823_/Y _3833_/X vssd1 vssd1 vccd1 vccd1 _3847_/A sky130_fd_sc_hd__o21ai_1
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3765_ _3752_/X _3757_/X _3809_/A vssd1 vssd1 vccd1 vccd1 _3778_/A sky130_fd_sc_hd__o21ai_2
X_5504_ _5504_/A _5525_/B _5504_/C vssd1 vssd1 vccd1 vccd1 _5509_/C sky130_fd_sc_hd__nand3_1
X_3696_ _3625_/Y _3691_/X _3695_/X vssd1 vssd1 vccd1 vccd1 _3696_/Y sky130_fd_sc_hd__a21oi_1
X_5435_ _5435_/A _5805_/B vssd1 vssd1 vccd1 vccd1 _5437_/A sky130_fd_sc_hd__nand2_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5366_ _5366_/A _5366_/B _5366_/C _5366_/D vssd1 vssd1 vccd1 vccd1 _5367_/B sky130_fd_sc_hd__nand4_1
X_5297_ _5297_/A _5297_/B _5297_/C vssd1 vssd1 vccd1 vccd1 _5297_/Y sky130_fd_sc_hd__nand3_2
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4317_ _4317_/A _4317_/B vssd1 vssd1 vccd1 vccd1 _4323_/A sky130_fd_sc_hd__nand2_1
X_4248_ _4110_/Y _4105_/B _4109_/Y vssd1 vssd1 vccd1 vccd1 _4250_/C sky130_fd_sc_hd__a21oi_2
X_4179_ _5553_/B vssd1 vssd1 vccd1 vccd1 _4179_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3550_ _4454_/B _4530_/A vssd1 vssd1 vccd1 vccd1 _3676_/A sky130_fd_sc_hd__nand2_2
X_5220_ _5833_/B _5810_/A _5411_/C _5833_/A vssd1 vssd1 vccd1 vccd1 _5220_/Y sky130_fd_sc_hd__a22oi_4
X_3481_ _3384_/X _3398_/X _3484_/A _3479_/Y _3480_/X vssd1 vssd1 vccd1 vccd1 _3482_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5151_ _5336_/A _5163_/B _5150_/Y vssd1 vssd1 vccd1 vccd1 _5151_/Y sky130_fd_sc_hd__a21oi_1
X_5082_ _5082_/A _5082_/B vssd1 vssd1 vccd1 vccd1 _5082_/Y sky130_fd_sc_hd__nand2_1
X_4102_ _4936_/A _5026_/A vssd1 vssd1 vccd1 vccd1 _4103_/B sky130_fd_sc_hd__nand2_2
X_4033_ _4029_/Y _4032_/Y _3964_/B vssd1 vssd1 vccd1 vccd1 _4177_/C sky130_fd_sc_hd__o21ai_2
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5984_ _5984_/A _5984_/B vssd1 vssd1 vccd1 vccd1 _5984_/X sky130_fd_sc_hd__or2_1
XFILLER_52_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4935_ _4935_/A _4935_/B _4935_/C _5119_/D vssd1 vssd1 vccd1 vccd1 _4935_/Y sky130_fd_sc_hd__nand4_4
XANTENNA_11 _6163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _6060_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4866_ _4731_/A _4860_/X _4745_/A vssd1 vssd1 vccd1 vccd1 _4866_/X sky130_fd_sc_hd__o21a_1
X_3817_ _3822_/A _3822_/B vssd1 vssd1 vccd1 vccd1 _3817_/Y sky130_fd_sc_hd__nand2_1
X_4797_ _4802_/B _4801_/B _4801_/A vssd1 vssd1 vccd1 vccd1 _4797_/Y sky130_fd_sc_hd__nand3_2
X_3748_ _4252_/A vssd1 vssd1 vccd1 vccd1 _4065_/A sky130_fd_sc_hd__buf_2
XFILLER_20_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3679_ _4873_/A _3711_/A vssd1 vssd1 vccd1 vccd1 _3679_/Y sky130_fd_sc_hd__nand2_2
X_5418_ _5430_/A _5614_/A _5429_/B vssd1 vssd1 vccd1 vccd1 _5418_/Y sky130_fd_sc_hd__a21oi_1
X_5349_ _5141_/C _6255_/B _5007_/A _5348_/X vssd1 vssd1 vccd1 vccd1 _5364_/B sky130_fd_sc_hd__a31oi_4
XFILLER_87_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4720_ _4712_/Y _4988_/B _4719_/Y vssd1 vssd1 vccd1 vccd1 _4720_/Y sky130_fd_sc_hd__a21oi_1
X_4651_ _4649_/Y _4650_/Y _4645_/Y _4817_/B _4806_/A vssd1 vssd1 vccd1 vccd1 _4652_/C
+ sky130_fd_sc_hd__o2111ai_1
Xinput31 b[6] vssd1 vssd1 vccd1 vccd1 _3536_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3602_ _6294_/B _3600_/C _3601_/A vssd1 vssd1 vccd1 vccd1 _3745_/A sky130_fd_sc_hd__a21oi_4
Xinput20 b[13] vssd1 vssd1 vccd1 vccd1 _4275_/A sky130_fd_sc_hd__clkbuf_1
X_4582_ _4579_/Y _4581_/Y _4573_/A vssd1 vssd1 vccd1 vccd1 _4586_/A sky130_fd_sc_hd__o21ai_1
X_3533_ _3533_/A _3533_/B _4931_/A _4229_/B vssd1 vssd1 vccd1 vccd1 _3657_/B sky130_fd_sc_hd__nand4_2
X_6252_ _6252_/A _6258_/A _6240_/X vssd1 vssd1 vccd1 vccd1 _6266_/C sky130_fd_sc_hd__or3b_1
X_3464_ _3574_/A _3574_/B _3574_/C vssd1 vssd1 vccd1 vccd1 _3486_/A sky130_fd_sc_hd__nand3_2
X_5203_ _5203_/A _5203_/B vssd1 vssd1 vccd1 vccd1 _5277_/A sky130_fd_sc_hd__nand2_1
X_6183_ _6183_/A _6183_/B _6182_/X vssd1 vssd1 vccd1 vccd1 _6222_/A sky130_fd_sc_hd__nor3b_4
X_3395_ _3315_/A _3315_/C _3394_/D _3597_/B vssd1 vssd1 vccd1 vccd1 _3395_/X sky130_fd_sc_hd__a2bb2o_1
X_5134_ _5134_/A _5134_/B vssd1 vssd1 vccd1 vccd1 _5141_/A sky130_fd_sc_hd__nand2_2
XFILLER_84_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5065_ _5065_/A _5065_/B vssd1 vssd1 vccd1 vccd1 _5067_/A sky130_fd_sc_hd__nand2_1
X_4016_ _6016_/A vssd1 vssd1 vccd1 vccd1 _6203_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5967_ _6255_/A vssd1 vssd1 vccd1 vccd1 _5967_/X sky130_fd_sc_hd__buf_2
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4918_ _4918_/A vssd1 vssd1 vccd1 vccd1 _5100_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5898_ _5872_/B _5872_/C _5872_/A vssd1 vssd1 vccd1 vccd1 _5898_/Y sky130_fd_sc_hd__a21oi_1
X_4849_ _4849_/A vssd1 vssd1 vccd1 vccd1 _4849_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ _4019_/A vssd1 vssd1 vccd1 vccd1 _3555_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_78_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5821_ _5821_/A vssd1 vssd1 vccd1 vccd1 _5957_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5752_ _5748_/X _5749_/Y _5751_/Y vssd1 vssd1 vccd1 vccd1 _5752_/X sky130_fd_sc_hd__o21a_1
XFILLER_22_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4703_ _4703_/A vssd1 vssd1 vccd1 vccd1 _4703_/X sky130_fd_sc_hd__buf_2
X_5683_ _5858_/C _6233_/C _6205_/B _5845_/A vssd1 vssd1 vccd1 vccd1 _5684_/B sky130_fd_sc_hd__a22oi_4
X_4634_ _4635_/A _4635_/B _4635_/C vssd1 vssd1 vccd1 vccd1 _4634_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4565_ _4564_/X _4561_/X _4554_/Y _4817_/A vssd1 vssd1 vccd1 vccd1 _4817_/B sky130_fd_sc_hd__o211ai_4
XFILLER_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3516_ _3509_/B _3516_/B _3516_/C vssd1 vssd1 vccd1 vccd1 _3522_/A sky130_fd_sc_hd__nand3b_2
X_4496_ _4648_/A _4498_/C _4647_/A vssd1 vssd1 vccd1 vccd1 _4499_/A sky130_fd_sc_hd__a21o_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6235_ _6235_/A _6235_/B _6235_/C _6235_/D vssd1 vssd1 vccd1 vccd1 _6235_/Y sky130_fd_sc_hd__nor4_4
X_3447_ _3348_/A _3358_/D _3347_/Y vssd1 vssd1 vccd1 vccd1 _3452_/A sky130_fd_sc_hd__a21oi_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6132_/C _6203_/D _6205_/B _6165_/A vssd1 vssd1 vccd1 vccd1 _6166_/Y sky130_fd_sc_hd__a22oi_2
X_3378_ _3398_/A _3398_/B _3398_/C vssd1 vssd1 vccd1 vccd1 _3483_/A sky130_fd_sc_hd__nand3_2
X_6097_ _6097_/A _6149_/B _6097_/C vssd1 vssd1 vccd1 vccd1 _6151_/A sky130_fd_sc_hd__nand3_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _5117_/A vssd1 vssd1 vccd1 vccd1 _5157_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5048_ _5048_/A _5053_/A _5237_/A _5240_/D vssd1 vssd1 vccd1 vccd1 _5081_/B sky130_fd_sc_hd__nand4_4
XFILLER_84_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4350_ _4194_/Y _4198_/Y _4219_/B vssd1 vssd1 vccd1 vccd1 _4399_/B sky130_fd_sc_hd__o21a_1
X_3301_ _3306_/A _3306_/B _3300_/C _3300_/D vssd1 vssd1 vccd1 vccd1 _3302_/C sky130_fd_sc_hd__a22o_1
X_4281_ _4298_/A _4298_/B _4298_/C _4298_/D vssd1 vssd1 vccd1 vccd1 _4281_/X sky130_fd_sc_hd__and4_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6020_ _6020_/A _6110_/A _6020_/C _6137_/B vssd1 vssd1 vccd1 vccd1 _6110_/B sky130_fd_sc_hd__nand4_2
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _4877_/B vssd1 vssd1 vccd1 vccd1 _5065_/A sky130_fd_sc_hd__clkbuf_2
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _3803_/A vssd1 vssd1 vccd1 vccd1 _3791_/C sky130_fd_sc_hd__buf_2
XFILLER_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5804_ _5810_/A vssd1 vssd1 vccd1 vccd1 _6020_/C sky130_fd_sc_hd__buf_2
XFILLER_62_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3996_ _3999_/A _3996_/B _3996_/C _3996_/D vssd1 vssd1 vccd1 vccd1 _4163_/C sky130_fd_sc_hd__nand4_2
X_5735_ _5588_/A _5588_/B _5588_/C vssd1 vssd1 vccd1 vccd1 _5735_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5666_ _5666_/A vssd1 vssd1 vccd1 vccd1 _5852_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4617_ _5026_/A _4777_/C vssd1 vssd1 vccd1 vccd1 _4618_/B sky130_fd_sc_hd__nand2_1
X_5597_ _5597_/A _5677_/A vssd1 vssd1 vccd1 vccd1 _5598_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4548_ _4365_/B _4533_/X _4547_/X _4529_/Y vssd1 vssd1 vccd1 vccd1 _4548_/X sky130_fd_sc_hd__o211a_1
X_4479_ _4489_/C _4641_/B _4468_/A vssd1 vssd1 vccd1 vccd1 _4479_/X sky130_fd_sc_hd__a21o_1
XFILLER_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6218_ _6218_/A _6218_/B vssd1 vssd1 vccd1 vccd1 _6218_/Y sky130_fd_sc_hd__xnor2_4
X_6149_ _6149_/A _6149_/B vssd1 vssd1 vccd1 vccd1 _6149_/Y sky130_fd_sc_hd__nand2_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3850_ _3840_/X _3996_/B _3849_/Y vssd1 vssd1 vccd1 vccd1 _3998_/C sky130_fd_sc_hd__o21ai_1
X_3781_ _3752_/X _3757_/X _3809_/A _3780_/X vssd1 vssd1 vccd1 vccd1 _3819_/C sky130_fd_sc_hd__o211ai_2
X_5520_ _5520_/A _5520_/B vssd1 vssd1 vccd1 vccd1 _5520_/X sky130_fd_sc_hd__and2_1
X_5451_ _5451_/A _5451_/B _5451_/C vssd1 vssd1 vccd1 vccd1 _5468_/C sky130_fd_sc_hd__nand3_2
X_4402_ _4945_/A _5037_/A vssd1 vssd1 vccd1 vccd1 _4402_/Y sky130_fd_sc_hd__nand2_1
X_5382_ _5603_/C _5677_/A _5382_/C vssd1 vssd1 vccd1 vccd1 _5383_/C sky130_fd_sc_hd__and3_1
X_4333_ _4333_/A _4333_/B _4333_/C vssd1 vssd1 vccd1 vccd1 _4334_/C sky130_fd_sc_hd__nand3_1
X_4264_ _4275_/A vssd1 vssd1 vccd1 vccd1 _4873_/B sky130_fd_sc_hd__buf_2
X_3215_ _3215_/A _3215_/B vssd1 vssd1 vccd1 vccd1 _3229_/A sky130_fd_sc_hd__nand2_1
X_6003_ _6125_/A _6003_/B vssd1 vssd1 vccd1 vccd1 _6004_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4195_ _5448_/A vssd1 vssd1 vccd1 vccd1 _6009_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3146_ _4355_/B vssd1 vssd1 vccd1 vccd1 _4186_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5718_ _5718_/A vssd1 vssd1 vccd1 vccd1 _6137_/B sky130_fd_sc_hd__buf_2
X_3979_ _3795_/Y _3791_/B _3879_/Y vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__a21oi_1
XFILLER_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5649_ _5622_/A _5622_/B _5622_/C _5629_/A vssd1 vssd1 vccd1 vccd1 _5649_/X sky130_fd_sc_hd__a31o_1
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput7 a[1] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4951_ _4951_/A _4951_/B vssd1 vssd1 vccd1 vccd1 _4951_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3902_ _3902_/A _3902_/B vssd1 vssd1 vccd1 vccd1 _3918_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4882_ _4885_/B _4885_/C _5594_/A _5411_/C vssd1 vssd1 vccd1 vccd1 _4882_/X sky130_fd_sc_hd__and4_1
X_3833_ _3993_/A _3833_/B vssd1 vssd1 vccd1 vccd1 _3833_/X sky130_fd_sc_hd__or2_1
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3764_ _3764_/A vssd1 vssd1 vccd1 vccd1 _3809_/A sky130_fd_sc_hd__clkbuf_2
X_5503_ _5502_/A _5494_/A _5502_/C vssd1 vssd1 vccd1 vccd1 _5504_/C sky130_fd_sc_hd__a21o_1
X_3695_ _4042_/B _3641_/A _6096_/C _3639_/X vssd1 vssd1 vccd1 vccd1 _3695_/X sky130_fd_sc_hd__a31o_1
X_5434_ _5436_/A _5435_/A _5436_/B _5434_/D vssd1 vssd1 vccd1 vccd1 _5464_/A sky130_fd_sc_hd__nand4_1
X_5365_ _5366_/A _5366_/B _5366_/C _5366_/D vssd1 vssd1 vccd1 vccd1 _5367_/A sky130_fd_sc_hd__a22o_1
X_5296_ _5296_/A _5925_/A _5436_/A _5296_/D vssd1 vssd1 vccd1 vccd1 _5297_/C sky130_fd_sc_hd__nand4_2
X_4316_ _4142_/Y _4144_/X _4123_/Y _4125_/Y vssd1 vssd1 vccd1 vccd1 _4317_/B sky130_fd_sc_hd__o22ai_1
X_4247_ _4247_/A vssd1 vssd1 vccd1 vccd1 _4302_/D sky130_fd_sc_hd__clkbuf_2
X_4178_ _4201_/C _4048_/C _4177_/X vssd1 vssd1 vccd1 vccd1 _4313_/A sky130_fd_sc_hd__a21oi_4
XFILLER_67_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3480_ _3486_/A _3486_/B _3479_/A vssd1 vssd1 vccd1 vccd1 _3480_/X sky130_fd_sc_hd__a21o_1
X_5150_ _4960_/Y _4938_/Y _4948_/Y vssd1 vssd1 vccd1 vccd1 _5150_/Y sky130_fd_sc_hd__o21ai_2
X_4101_ _4096_/X _4098_/Y _4130_/A _4100_/X vssd1 vssd1 vccd1 vccd1 _4124_/A sky130_fd_sc_hd__o22ai_4
X_5081_ _5081_/A _5081_/B _5087_/C _5372_/C vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__and4_1
X_4032_ _4540_/A _5792_/A _5794_/B _3960_/B vssd1 vssd1 vccd1 vccd1 _4032_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5983_ _5984_/A _5984_/B vssd1 vssd1 vccd1 vccd1 _5983_/Y sky130_fd_sc_hd__nand2_1
X_4934_ _4417_/X _5453_/B _4928_/X _5124_/A _4933_/X vssd1 vssd1 vccd1 vccd1 _4934_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA_12 _3171_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _6118_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4865_ _5088_/A _5088_/B _4865_/C vssd1 vssd1 vccd1 vccd1 _4865_/Y sky130_fd_sc_hd__nand3_2
X_3816_ _3809_/Y _3810_/Y _3811_/Y _3815_/Y vssd1 vssd1 vccd1 vccd1 _3822_/B sky130_fd_sc_hd__o211ai_4
X_4796_ _4796_/A _4796_/B vssd1 vssd1 vccd1 vccd1 _4802_/B sky130_fd_sc_hd__nor2_1
X_3747_ _3747_/A _3747_/B vssd1 vssd1 vccd1 vccd1 _3755_/A sky130_fd_sc_hd__nand2_1
X_3678_ _4939_/A _5263_/C _3676_/Y _3677_/Y vssd1 vssd1 vccd1 vccd1 _3684_/A sky130_fd_sc_hd__a22oi_4
X_5417_ _5614_/B _5614_/C vssd1 vssd1 vccd1 vccd1 _5429_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5348_ _5511_/C _5465_/C _5506_/A _5348_/D vssd1 vssd1 vccd1 vccd1 _5348_/X sky130_fd_sc_hd__and4_1
X_5279_ _5221_/X _5226_/X _5274_/Y _5275_/Y vssd1 vssd1 vccd1 vccd1 _5485_/B sky130_fd_sc_hd__o22ai_2
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4650_ _4466_/C _4640_/Y _4641_/Y _4639_/B vssd1 vssd1 vccd1 vccd1 _4650_/Y sky130_fd_sc_hd__o211ai_4
Xinput10 a[4] vssd1 vssd1 vccd1 vccd1 _3897_/A sky130_fd_sc_hd__clkbuf_4
X_3601_ _3601_/A _3601_/B vssd1 vssd1 vccd1 vccd1 _3601_/Y sky130_fd_sc_hd__xnor2_1
Xinput21 b[14] vssd1 vssd1 vccd1 vccd1 _4569_/A sky130_fd_sc_hd__clkbuf_2
Xinput32 b[7] vssd1 vssd1 vccd1 vccd1 _3766_/A sky130_fd_sc_hd__buf_4
X_4581_ _4581_/A _4731_/A vssd1 vssd1 vccd1 vccd1 _4581_/Y sky130_fd_sc_hd__nor2_1
X_3532_ _3758_/B vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__clkbuf_2
X_6251_ _6251_/A _6251_/B vssd1 vssd1 vccd1 vccd1 _6251_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3463_ _3459_/Y _3462_/Y _3446_/X _3465_/A _3465_/B vssd1 vssd1 vccd1 vccd1 _3574_/C
+ sky130_fd_sc_hd__o2111ai_4
X_6182_ _6149_/Y _6181_/X _6151_/Y vssd1 vssd1 vccd1 vccd1 _6182_/X sky130_fd_sc_hd__a21o_1
X_5202_ _5202_/A _5202_/B vssd1 vssd1 vccd1 vccd1 _5203_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3394_ _3315_/A _3394_/B _3394_/C _3394_/D vssd1 vssd1 vccd1 vccd1 _3597_/A sky130_fd_sc_hd__nand4b_2
X_5133_ _4936_/A input4/X input5/X _3867_/A vssd1 vssd1 vccd1 vccd1 _5136_/A sky130_fd_sc_hd__a22o_1
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5064_ _5064_/A _5211_/B vssd1 vssd1 vccd1 vccd1 _5070_/A sky130_fd_sc_hd__nand2_2
X_4015_ _5810_/B vssd1 vssd1 vccd1 vccd1 _6016_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ _5966_/A _5966_/B _5966_/C vssd1 vssd1 vccd1 vccd1 _5969_/B sky130_fd_sc_hd__nand3_1
X_5897_ _5897_/A _5897_/B vssd1 vssd1 vccd1 vccd1 _5897_/Y sky130_fd_sc_hd__xnor2_4
X_4917_ _4917_/A _4917_/B _4917_/C vssd1 vssd1 vccd1 vccd1 _5100_/A sky130_fd_sc_hd__nand3_2
X_4848_ _4848_/A _4848_/B vssd1 vssd1 vccd1 vccd1 _4849_/A sky130_fd_sc_hd__and2_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4779_ _5530_/A _4779_/B vssd1 vssd1 vccd1 vccd1 _4779_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5820_ _5865_/B _5865_/C vssd1 vssd1 vccd1 vccd1 _5821_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5751_ _5556_/Y _5694_/X _5750_/Y vssd1 vssd1 vccd1 vccd1 _5751_/Y sky130_fd_sc_hd__o21ai_2
X_4702_ _4702_/A _4702_/B _4702_/C vssd1 vssd1 vccd1 vccd1 _4722_/A sky130_fd_sc_hd__nand3_4
X_5682_ _6165_/D vssd1 vssd1 vccd1 vccd1 _6205_/B sky130_fd_sc_hd__clkbuf_4
X_4633_ _4417_/X _3797_/X _4405_/Y _4618_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4635_/C
+ sky130_fd_sc_hd__o32a_2
X_4564_ _4564_/A _4564_/B _4564_/C vssd1 vssd1 vccd1 vccd1 _4564_/X sky130_fd_sc_hd__and3_2
X_3515_ _3508_/D _3641_/A _3514_/Y vssd1 vssd1 vccd1 vccd1 _3516_/C sky130_fd_sc_hd__a21o_1
X_6234_ _6235_/A _6235_/B _6235_/C _6235_/D vssd1 vssd1 vccd1 vccd1 _6234_/X sky130_fd_sc_hd__o22a_1
X_4495_ _4495_/A _4495_/B vssd1 vssd1 vccd1 vccd1 _4647_/A sky130_fd_sc_hd__nand2_2
X_3446_ _3446_/A vssd1 vssd1 vccd1 vccd1 _3446_/X sky130_fd_sc_hd__clkbuf_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6165_ _6165_/A _6165_/B _6203_/D _6165_/D vssd1 vssd1 vccd1 vccd1 _6165_/X sky130_fd_sc_hd__and4_1
X_3377_ _3362_/Y _3367_/Y _3370_/X _3477_/A _3376_/Y vssd1 vssd1 vccd1 vccd1 _3398_/C
+ sky130_fd_sc_hd__o2111ai_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _5116_/A _5116_/B _5116_/C vssd1 vssd1 vccd1 vccd1 _5117_/A sky130_fd_sc_hd__nand3_1
X_6096_ _6096_/A _6253_/A _6096_/C vssd1 vssd1 vccd1 vccd1 _6097_/C sky130_fd_sc_hd__and3_2
X_5047_ _5238_/A vssd1 vssd1 vccd1 vccd1 _5240_/D sky130_fd_sc_hd__buf_2
XFILLER_72_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5949_ _5949_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5952_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3300_ _3306_/A _3306_/B _3300_/C _3300_/D vssd1 vssd1 vccd1 vccd1 _3302_/B sky130_fd_sc_hd__nand4_1
X_4280_ _4294_/B vssd1 vssd1 vccd1 vccd1 _4298_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _3897_/A vssd1 vssd1 vccd1 vccd1 _4877_/B sky130_fd_sc_hd__clkbuf_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _4714_/A vssd1 vssd1 vccd1 vccd1 _3803_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5803_ _5816_/B _5945_/A vssd1 vssd1 vccd1 vccd1 _5814_/A sky130_fd_sc_hd__nand2_1
X_3995_ _3999_/A _3996_/B _3996_/C _3996_/D vssd1 vssd1 vccd1 vccd1 _4166_/A sky130_fd_sc_hd__a22oi_2
XFILLER_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5734_ _5728_/A _5728_/B _5733_/Y vssd1 vssd1 vccd1 vccd1 _5734_/Y sky130_fd_sc_hd__a21oi_2
X_5665_ _5657_/Y _5659_/Y _5661_/Y _5664_/X vssd1 vssd1 vccd1 vccd1 _5673_/B sky130_fd_sc_hd__o211ai_4
X_4616_ _4935_/A _5211_/A vssd1 vssd1 vccd1 vccd1 _4618_/A sky130_fd_sc_hd__nand2_1
X_5596_ _5596_/A _5596_/B _5676_/A _5681_/A vssd1 vssd1 vccd1 vccd1 _5604_/B sky130_fd_sc_hd__nand4_2
X_4547_ _4547_/A _5704_/B vssd1 vssd1 vccd1 vccd1 _4547_/X sky130_fd_sc_hd__and2_1
X_4478_ _4478_/A _4640_/A _4640_/B vssd1 vssd1 vccd1 vccd1 _4489_/C sky130_fd_sc_hd__nand3_1
X_6217_ _6224_/A _6197_/B _6190_/X vssd1 vssd1 vccd1 vccd1 _6218_/B sky130_fd_sc_hd__o21ai_2
X_3429_ _4571_/B _4228_/A vssd1 vssd1 vccd1 vccd1 _3429_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6148_ _6148_/A _6148_/B vssd1 vssd1 vccd1 vccd1 _6151_/B sky130_fd_sc_hd__nand2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6079_ _6079_/A _6137_/B vssd1 vssd1 vccd1 vccd1 _6084_/A sky130_fd_sc_hd__nand2_1
XFILLER_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3780_ _3768_/Y _3771_/X _3776_/Y vssd1 vssd1 vccd1 vccd1 _3780_/X sky130_fd_sc_hd__o21a_2
X_5450_ _5291_/X _5542_/A _5712_/A _6010_/A _5445_/Y vssd1 vssd1 vccd1 vccd1 _5451_/C
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4401_ _5397_/A _5119_/A vssd1 vssd1 vccd1 vccd1 _4411_/B sky130_fd_sc_hd__nand2_1
X_5381_ _5246_/X _5598_/A _5263_/C _6001_/C _5375_/Y vssd1 vssd1 vccd1 vccd1 _5383_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4332_ _4043_/C _4043_/A _4043_/B _4054_/X vssd1 vssd1 vccd1 vccd1 _4333_/C sky130_fd_sc_hd__a31o_1
X_4263_ _4861_/A _5207_/B vssd1 vssd1 vccd1 vccd1 _4429_/A sky130_fd_sc_hd__nand2_2
X_6002_ _6124_/A _6002_/B vssd1 vssd1 vccd1 vccd1 _6004_/A sky130_fd_sc_hd__nand2_1
X_3214_ _4067_/A _4708_/B vssd1 vssd1 vccd1 vccd1 _3215_/B sky130_fd_sc_hd__nand2_2
X_4194_ _4197_/B _4182_/Y _4197_/A vssd1 vssd1 vccd1 vccd1 _4194_/Y sky130_fd_sc_hd__a21oi_4
X_3145_ _3473_/A vssd1 vssd1 vccd1 vccd1 _4355_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ _3973_/A _3973_/B _3975_/B vssd1 vssd1 vccd1 vccd1 _3990_/A sky130_fd_sc_hd__a21o_1
X_5717_ _5719_/C _5933_/D _5719_/D _5719_/A vssd1 vssd1 vccd1 vccd1 _5733_/A sky130_fd_sc_hd__a22o_1
X_5648_ _5638_/A _5640_/D _5647_/Y vssd1 vssd1 vccd1 vccd1 _5773_/A sky130_fd_sc_hd__a21o_1
X_5579_ _5674_/A _5674_/B _5654_/A _5585_/A vssd1 vssd1 vccd1 vccd1 _5584_/B sky130_fd_sc_hd__o211ai_4
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput8 a[2] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4950_ _4950_/A _4950_/B vssd1 vssd1 vccd1 vccd1 _4951_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3901_ _3902_/A _3902_/B _3918_/A vssd1 vssd1 vccd1 vccd1 _3901_/X sky130_fd_sc_hd__a21o_1
XFILLER_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4881_ _5541_/B vssd1 vssd1 vccd1 vccd1 _5411_/C sky130_fd_sc_hd__clkbuf_4
X_3832_ _3829_/X _3830_/Y _3691_/X _3824_/Y vssd1 vssd1 vccd1 vccd1 _3833_/B sky130_fd_sc_hd__o211a_1
X_5502_ _5502_/A _5525_/A _5502_/C vssd1 vssd1 vccd1 vccd1 _5525_/B sky130_fd_sc_hd__nand3_1
X_3763_ _3759_/Y _3760_/Y _3761_/Y _3762_/X vssd1 vssd1 vccd1 vccd1 _3764_/A sky130_fd_sc_hd__o211ai_4
X_3694_ _5994_/B vssd1 vssd1 vccd1 vccd1 _6096_/C sky130_fd_sc_hd__buf_2
X_5433_ _5218_/A _5218_/B _5218_/C _5281_/C vssd1 vssd1 vccd1 vccd1 _5433_/Y sky130_fd_sc_hd__a31oi_2
X_5364_ _5364_/A _5364_/B vssd1 vssd1 vccd1 vccd1 _5513_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4315_ _4315_/A _4315_/B _4315_/C vssd1 vssd1 vccd1 vccd1 _4333_/A sky130_fd_sc_hd__nand3_2
X_5295_ _5296_/D _5296_/A _4255_/Y _5446_/A vssd1 vssd1 vccd1 vccd1 _5297_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4246_ _4232_/Y _4243_/X _4244_/Y _4245_/Y vssd1 vssd1 vccd1 vccd1 _4247_/A sky130_fd_sc_hd__o211ai_4
X_4177_ _4177_/A _4177_/B _4177_/C vssd1 vssd1 vccd1 vccd1 _4177_/X sky130_fd_sc_hd__and3_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5080_ _5080_/A _5080_/B _5248_/A _5794_/C vssd1 vssd1 vccd1 vccd1 _5080_/X sky130_fd_sc_hd__and4_1
X_4100_ _4100_/A _4100_/B _4100_/C vssd1 vssd1 vccd1 vccd1 _4100_/X sky130_fd_sc_hd__and3_1
XFILLER_84_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4031_ _5448_/A vssd1 vssd1 vccd1 vccd1 _5794_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5982_ _6193_/A _5982_/B vssd1 vssd1 vccd1 vccd1 _5982_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4933_ _4933_/A vssd1 vssd1 vccd1 vccd1 _4933_/X sky130_fd_sc_hd__buf_2
XFILLER_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_13 _6273_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4864_ _4860_/X _5258_/A _4277_/C _5575_/B _5087_/A vssd1 vssd1 vccd1 vccd1 _4865_/C
+ sky130_fd_sc_hd__o2111ai_1
XANTENNA_24 _3245_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3815_ _3813_/Y _3814_/X _3778_/A vssd1 vssd1 vccd1 vccd1 _3815_/Y sky130_fd_sc_hd__o21ai_1
X_4795_ _4795_/A _4795_/B vssd1 vssd1 vccd1 vccd1 _4795_/Y sky130_fd_sc_hd__nand2_2
X_3746_ input1/X _4252_/A vssd1 vssd1 vccd1 vccd1 _3747_/B sky130_fd_sc_hd__nand2_2
XFILLER_21_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5416_ _5411_/X _5213_/X _5414_/Y _5415_/X vssd1 vssd1 vccd1 vccd1 _5614_/C sky130_fd_sc_hd__o22ai_4
X_3677_ _3677_/A _5372_/B _4363_/B _5132_/B vssd1 vssd1 vccd1 vccd1 _3677_/Y sky130_fd_sc_hd__nand4_2
X_5347_ _5347_/A vssd1 vssd1 vccd1 vccd1 _5465_/C sky130_fd_sc_hd__clkbuf_2
X_5278_ _5278_/A _5278_/B vssd1 vssd1 vccd1 vccd1 _5485_/A sky130_fd_sc_hd__nand2_1
X_4229_ _5397_/A _4229_/B vssd1 vssd1 vccd1 vccd1 _4239_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput11 a[5] vssd1 vssd1 vccd1 vccd1 _3322_/A sky130_fd_sc_hd__clkbuf_4
Xinput22 b[15] vssd1 vssd1 vccd1 vccd1 _4578_/A sky130_fd_sc_hd__buf_4
X_3600_ _6294_/A _6294_/B _3600_/C vssd1 vssd1 vccd1 vccd1 _3601_/B sky130_fd_sc_hd__nand3_1
X_4580_ _4855_/B _4863_/A vssd1 vssd1 vccd1 vccd1 _4731_/A sky130_fd_sc_hd__nand2_2
Xinput33 b[8] vssd1 vssd1 vccd1 vccd1 _3903_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3531_ _3658_/A vssd1 vssd1 vccd1 vccd1 _3564_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6250_ _6224_/B _6223_/X _6274_/A _6197_/B _6275_/C vssd1 vssd1 vccd1 vccd1 _6251_/B
+ sky130_fd_sc_hd__o221a_1
X_3462_ _3461_/Y _3439_/A _3452_/A vssd1 vssd1 vccd1 vccd1 _3462_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6181_ _6097_/A _6149_/B _6097_/C _6148_/A _6148_/B vssd1 vssd1 vccd1 vccd1 _6181_/X
+ sky130_fd_sc_hd__a32o_1
X_5201_ _5200_/Y _5117_/A _5107_/A vssd1 vssd1 vccd1 vccd1 _5323_/A sky130_fd_sc_hd__a21boi_1
X_3393_ _3315_/A _3598_/B _3394_/D _3597_/B vssd1 vssd1 vccd1 vccd1 _3598_/C sky130_fd_sc_hd__a2bb2oi_2
X_5132_ _5132_/A _5132_/B _5532_/C _5532_/D vssd1 vssd1 vccd1 vccd1 _5141_/B sky130_fd_sc_hd__nand4_4
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5063_ _5207_/B vssd1 vssd1 vccd1 vccd1 _5211_/B sky130_fd_sc_hd__clkbuf_2
X_4014_ _5299_/C vssd1 vssd1 vccd1 vccd1 _5810_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_92_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5965_ _5956_/A _5956_/B _5964_/Y vssd1 vssd1 vccd1 vccd1 _5966_/B sky130_fd_sc_hd__o21ai_1
XFILLER_25_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5896_ _5974_/B _5780_/B _5974_/A vssd1 vssd1 vccd1 vccd1 _5897_/B sky130_fd_sc_hd__a21bo_1
X_4916_ _4916_/A _5534_/A _5578_/A vssd1 vssd1 vccd1 vccd1 _4917_/C sky130_fd_sc_hd__nand3_2
X_4847_ _5518_/A _4847_/B vssd1 vssd1 vccd1 vccd1 _4848_/B sky130_fd_sc_hd__or2_1
XFILLER_33_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4778_ _4255_/Y _3634_/A _4784_/A _4784_/B vssd1 vssd1 vccd1 vccd1 _4781_/B sky130_fd_sc_hd__o211ai_2
X_3729_ _3730_/A _3730_/B _3729_/C vssd1 vssd1 vccd1 vccd1 _3732_/A sky130_fd_sc_hd__and3_1
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5750_ _5734_/Y _5738_/Y _5723_/Y vssd1 vssd1 vccd1 vccd1 _5750_/Y sky130_fd_sc_hd__o21ai_1
X_4701_ _4703_/A _4698_/Y _4700_/Y vssd1 vssd1 vccd1 vccd1 _4702_/C sky130_fd_sc_hd__o21bai_1
X_5681_ _5681_/A vssd1 vssd1 vccd1 vccd1 _6165_/D sky130_fd_sc_hd__clkbuf_2
X_4632_ _4632_/A _4795_/A vssd1 vssd1 vccd1 vccd1 _4639_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4563_ _4554_/Y _4817_/A _4562_/X vssd1 vssd1 vccd1 vccd1 _4806_/A sky130_fd_sc_hd__a21o_1
X_4494_ _4494_/A _4494_/B _4494_/C vssd1 vssd1 vccd1 vccd1 _4502_/A sky130_fd_sc_hd__nand3_4
X_3514_ _3514_/A _5578_/A vssd1 vssd1 vccd1 vccd1 _3514_/Y sky130_fd_sc_hd__nand2_1
X_6233_ _6233_/A _6233_/B _6233_/C _6253_/A vssd1 vssd1 vccd1 vccd1 _6235_/D sky130_fd_sc_hd__and4_2
X_3445_ _3445_/A _3445_/B _3445_/C vssd1 vssd1 vccd1 vccd1 _3446_/A sky130_fd_sc_hd__nand3_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6164_/A _6164_/B vssd1 vssd1 vccd1 vccd1 _6180_/C sky130_fd_sc_hd__nand2_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3440_/B _3347_/Y _3374_/X _3375_/X vssd1 vssd1 vccd1 vccd1 _3376_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_84_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6205_/B vssd1 vssd1 vccd1 vccd1 _6253_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5115_ _4893_/C _5113_/Y _5114_/Y vssd1 vssd1 vccd1 vccd1 _5116_/C sky130_fd_sc_hd__o21ai_1
X_5046_ _5046_/A _5046_/B vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__nand2_2
XFILLER_84_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5948_ _5949_/A _5949_/B _5948_/C _5948_/D vssd1 vssd1 vccd1 vccd1 _5960_/B sky130_fd_sc_hd__nand4_2
XFILLER_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5879_ _5879_/A _5879_/B _5879_/C vssd1 vssd1 vccd1 vccd1 _5879_/Y sky130_fd_sc_hd__nand3_2
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3230_/A _3230_/B _3230_/C vssd1 vssd1 vccd1 vccd1 _3240_/B sky130_fd_sc_hd__nand3_2
XFILLER_94_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _3256_/A vssd1 vssd1 vccd1 vccd1 _4714_/A sky130_fd_sc_hd__buf_2
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5802_ _5802_/A vssd1 vssd1 vccd1 vccd1 _5945_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3994_ _3994_/A _4160_/C vssd1 vssd1 vccd1 vccd1 _3996_/D sky130_fd_sc_hd__nand2_1
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5733_ _5733_/A _5733_/B vssd1 vssd1 vccd1 vccd1 _5733_/Y sky130_fd_sc_hd__nand2_1
X_5664_ _5666_/A _5825_/B _5656_/Y vssd1 vssd1 vccd1 vccd1 _5664_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4615_ _5212_/A vssd1 vssd1 vccd1 vccd1 _5582_/A sky130_fd_sc_hd__clkbuf_4
X_5595_ _3310_/C _5678_/A _6124_/B _5681_/A _5604_/A vssd1 vssd1 vccd1 vccd1 _5595_/X
+ sky130_fd_sc_hd__a41o_1
X_4546_ _4689_/A _4689_/B vssd1 vssd1 vccd1 vccd1 _4546_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4477_ _4463_/A _4463_/B _4474_/Y _4476_/X vssd1 vssd1 vccd1 vccd1 _4640_/B sky130_fd_sc_hd__o2bb2ai_1
X_6216_ _6222_/A _6222_/B _6215_/Y vssd1 vssd1 vccd1 vccd1 _6218_/A sky130_fd_sc_hd__o21ai_2
X_3428_ _3711_/A vssd1 vssd1 vccd1 vccd1 _4228_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6147_ _6097_/A _6149_/B _6097_/C _6148_/A _6148_/B vssd1 vssd1 vccd1 vccd1 _6147_/Y
+ sky130_fd_sc_hd__a32oi_2
X_3359_ _3359_/A _3359_/B _3359_/C vssd1 vssd1 vccd1 vccd1 _3360_/A sky130_fd_sc_hd__nand3_2
XFILLER_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6078_ _6078_/A _6078_/B vssd1 vssd1 vccd1 vccd1 _6081_/B sky130_fd_sc_hd__nand2_1
X_5029_ _5029_/A _5029_/B vssd1 vssd1 vccd1 vccd1 _5208_/A sky130_fd_sc_hd__nand2_4
XFILLER_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4400_ _4400_/A _4400_/B _4400_/C vssd1 vssd1 vccd1 vccd1 _4495_/B sky130_fd_sc_hd__nand3_2
X_5380_ _5919_/B vssd1 vssd1 vccd1 vccd1 _6001_/C sky130_fd_sc_hd__clkbuf_4
X_4331_ _4331_/A _4331_/B vssd1 vssd1 vccd1 vccd1 _4334_/B sky130_fd_sc_hd__nand2_1
X_4262_ _4275_/A vssd1 vssd1 vccd1 vccd1 _5207_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3213_ _3356_/A vssd1 vssd1 vccd1 vccd1 _4708_/B sky130_fd_sc_hd__clkbuf_4
X_6001_ _6125_/A _6124_/A _6001_/C _6003_/B vssd1 vssd1 vccd1 vccd1 _6006_/D sky130_fd_sc_hd__nand4_4
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4193_ _4193_/A _5925_/A vssd1 vssd1 vccd1 vccd1 _4197_/A sky130_fd_sc_hd__nand2_2
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3144_ _3179_/C vssd1 vssd1 vccd1 vccd1 _3190_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_67_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3977_ _3977_/A vssd1 vssd1 vccd1 vccd1 _4160_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5716_ _5724_/A _5728_/B _5729_/A _5729_/B vssd1 vssd1 vccd1 vccd1 _5748_/A sky130_fd_sc_hd__o2bb2ai_1
X_5647_ _5635_/B _5635_/C _5635_/A vssd1 vssd1 vccd1 vccd1 _5647_/Y sky130_fd_sc_hd__a21oi_1
X_5578_ _5578_/A _5688_/A vssd1 vssd1 vccd1 vccd1 _5585_/A sky130_fd_sc_hd__nand2_2
X_4529_ _4529_/A _4529_/B vssd1 vssd1 vccd1 vccd1 _4529_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput9 a[3] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_91_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3900_ _5064_/A _4228_/A vssd1 vssd1 vccd1 vccd1 _3918_/A sky130_fd_sc_hd__nand2_2
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4880_ _4880_/A vssd1 vssd1 vccd1 vccd1 _5594_/A sky130_fd_sc_hd__clkbuf_4
X_3831_ _3691_/X _3824_/Y _3829_/X _3830_/Y vssd1 vssd1 vccd1 vccd1 _3993_/A sky130_fd_sc_hd__a211oi_2
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3762_ _3755_/A _3755_/B _3758_/Y vssd1 vssd1 vccd1 vccd1 _3762_/X sky130_fd_sc_hd__a21o_1
X_5501_ _5337_/X _5335_/B _5340_/Y vssd1 vssd1 vccd1 vccd1 _5504_/A sky130_fd_sc_hd__a21o_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3693_ _5656_/A vssd1 vssd1 vccd1 vccd1 _5994_/B sky130_fd_sc_hd__buf_2
X_5432_ _5218_/A _5218_/B _5218_/C vssd1 vssd1 vccd1 vccd1 _5432_/Y sky130_fd_sc_hd__a21oi_4
X_5363_ _5363_/A _5363_/B vssd1 vssd1 vccd1 vccd1 _5363_/Y sky130_fd_sc_hd__xnor2_4
X_4314_ _4322_/A _4322_/B _4312_/Y _4313_/X vssd1 vssd1 vccd1 vccd1 _4315_/C sky130_fd_sc_hd__o2bb2ai_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5294_ _5120_/A _5128_/B _5121_/Y vssd1 vssd1 vccd1 vccd1 _5297_/A sky130_fd_sc_hd__a21oi_2
X_4245_ _4238_/Y _4240_/A _3448_/X _3634_/A vssd1 vssd1 vccd1 vccd1 _4245_/Y sky130_fd_sc_hd__o2bb2ai_1
X_4176_ _4176_/A _5299_/C vssd1 vssd1 vccd1 vccd1 _4201_/C sky130_fd_sc_hd__and2_1
XFILLER_27_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4030_ input2/X vssd1 vssd1 vccd1 vccd1 _5448_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5981_ _5981_/A _5981_/B vssd1 vssd1 vccd1 vccd1 _5982_/B sky130_fd_sc_hd__nand2_4
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4932_ _4932_/A _4932_/B vssd1 vssd1 vccd1 vccd1 _4933_/A sky130_fd_sc_hd__nand2_1
XFILLER_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_14 _3317_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4863_ _4863_/A vssd1 vssd1 vccd1 vccd1 _5575_/B sky130_fd_sc_hd__buf_4
XANTENNA_25 _6295_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3814_ _3814_/A _5678_/B _5511_/C vssd1 vssd1 vccd1 vccd1 _3814_/X sky130_fd_sc_hd__and3_1
X_4794_ _4794_/A _4794_/B vssd1 vssd1 vccd1 vccd1 _4794_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3745_ _3745_/A _3745_/B vssd1 vssd1 vccd1 vccd1 _3745_/X sky130_fd_sc_hd__xor2_4
XFILLER_9_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5415_ _3634_/X _5407_/Y _5408_/Y _5402_/Y vssd1 vssd1 vccd1 vccd1 _5415_/X sky130_fd_sc_hd__o211a_1
X_3676_ _3676_/A _3676_/B vssd1 vssd1 vccd1 vccd1 _3676_/Y sky130_fd_sc_hd__nand2_2
X_5346_ _5351_/A _5364_/A vssd1 vssd1 vccd1 vccd1 _5350_/A sky130_fd_sc_hd__nand2_1
X_5277_ _5277_/A _5277_/B _5277_/C vssd1 vssd1 vccd1 vccd1 _5277_/Y sky130_fd_sc_hd__nand3_2
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4228_ _4228_/A _5026_/B vssd1 vssd1 vccd1 vccd1 _4239_/A sky130_fd_sc_hd__nand2_1
XFILLER_68_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4159_ _4159_/A _4159_/B _4159_/C vssd1 vssd1 vccd1 vccd1 _4165_/A sky130_fd_sc_hd__nand3_1
XFILLER_46_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 a[6] vssd1 vssd1 vccd1 vccd1 _4901_/A sky130_fd_sc_hd__buf_4
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput23 b[16] vssd1 vssd1 vccd1 vccd1 _4732_/A sky130_fd_sc_hd__clkbuf_4
X_3530_ _3530_/A _3530_/B vssd1 vssd1 vccd1 vccd1 _3658_/A sky130_fd_sc_hd__nand2_1
Xinput34 b[9] vssd1 vssd1 vccd1 vccd1 _4407_/A sky130_fd_sc_hd__clkbuf_4
X_3461_ _5240_/B _4530_/A vssd1 vssd1 vccd1 vccd1 _3461_/Y sky130_fd_sc_hd__nand2_2
X_5200_ _5200_/A _5200_/B vssd1 vssd1 vccd1 vccd1 _5200_/Y sky130_fd_sc_hd__nand2_1
X_6180_ _6180_/A _6180_/B _6180_/C vssd1 vssd1 vccd1 vccd1 _6183_/B sky130_fd_sc_hd__and3_1
X_3392_ _3392_/A _3392_/B _3392_/C _3392_/D vssd1 vssd1 vccd1 vccd1 _3597_/B sky130_fd_sc_hd__nand4_4
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5131_ _5131_/A vssd1 vssd1 vccd1 vccd1 _5366_/A sky130_fd_sc_hd__buf_2
X_5062_ _5062_/A _5062_/B _5062_/C vssd1 vssd1 vccd1 vccd1 _5095_/B sky130_fd_sc_hd__nand3_4
XFILLER_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4013_ input4/X vssd1 vssd1 vccd1 vccd1 _5299_/C sky130_fd_sc_hd__buf_2
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5964_ _5956_/A _5956_/B _5962_/Y vssd1 vssd1 vccd1 vccd1 _5964_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_40_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5895_ _5974_/C _5974_/D vssd1 vssd1 vccd1 vccd1 _5897_/A sky130_fd_sc_hd__nand2_2
X_4915_ _4903_/A _4903_/B _4907_/X _4776_/B vssd1 vssd1 vccd1 vccd1 _4916_/A sky130_fd_sc_hd__o2bb2ai_1
XFILLER_33_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4846_ _4840_/X _4841_/X _4842_/Y _4523_/S vssd1 vssd1 vccd1 vccd1 _4847_/B sky130_fd_sc_hd__o22a_2
XFILLER_20_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4777_ _5026_/A _5026_/B _4777_/C _4777_/D vssd1 vssd1 vccd1 vccd1 _4784_/B sky130_fd_sc_hd__nand4_4
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3728_ _3731_/C _3829_/C vssd1 vssd1 vccd1 vccd1 _3729_/C sky130_fd_sc_hd__nand2_1
X_3659_ _3766_/A vssd1 vssd1 vccd1 vccd1 _3669_/A sky130_fd_sc_hd__inv_2
X_5329_ _5366_/C _5366_/D _5328_/A vssd1 vssd1 vccd1 vccd1 _5329_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5680_ _6065_/D vssd1 vssd1 vccd1 vccd1 _6233_/C sky130_fd_sc_hd__clkbuf_2
X_4700_ _4700_/A _5288_/B vssd1 vssd1 vccd1 vccd1 _4700_/Y sky130_fd_sc_hd__nand2_2
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4631_ _4631_/A _4631_/B vssd1 vssd1 vccd1 vccd1 _4795_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4562_ _4564_/C _4564_/A _4564_/B _4561_/X vssd1 vssd1 vccd1 vccd1 _4562_/X sky130_fd_sc_hd__a31o_2
XFILLER_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4493_ _4495_/A _4495_/B _4481_/A _4498_/C vssd1 vssd1 vccd1 vccd1 _4494_/C sky130_fd_sc_hd__a22o_1
X_3513_ _3186_/X _3512_/X _3508_/D _3641_/A vssd1 vssd1 vccd1 vccd1 _3516_/B sky130_fd_sc_hd__o211ai_1
X_6232_ _5348_/D _6255_/C _6253_/A _5506_/A vssd1 vssd1 vccd1 vccd1 _6235_/C sky130_fd_sc_hd__a22oi_4
X_3444_ _3441_/X _3448_/A _3342_/B _3530_/A _3443_/X vssd1 vssd1 vccd1 vccd1 _3445_/C
+ sky130_fd_sc_hd__o221ai_2
X_6163_ _6219_/A _6163_/B vssd1 vssd1 vccd1 vccd1 _6163_/X sky130_fd_sc_hd__xor2_4
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _3358_/D _3440_/A _3348_/A vssd1 vssd1 vccd1 vccd1 _3375_/X sky130_fd_sc_hd__a21o_1
X_6094_ _6094_/A _6094_/B _6149_/A vssd1 vssd1 vccd1 vccd1 _6149_/B sky130_fd_sc_hd__nand3_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5114_ _4919_/Y _4922_/X _4894_/A vssd1 vssd1 vccd1 vccd1 _5114_/Y sky130_fd_sc_hd__o21ai_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5045_ _5045_/A _5238_/A vssd1 vssd1 vccd1 vccd1 _5046_/B sky130_fd_sc_hd__nand2_2
XFILLER_38_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5947_ _5944_/A _5944_/B _5945_/A _5940_/Y _5943_/Y vssd1 vssd1 vccd1 vccd1 _5948_/D
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5878_ _5869_/Y _5877_/X _5866_/Y _5865_/X _5859_/Y vssd1 vssd1 vccd1 vccd1 _5879_/C
+ sky130_fd_sc_hd__o221ai_2
XFILLER_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4829_ _4829_/A vssd1 vssd1 vccd1 vccd1 _4830_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _3204_/B vssd1 vssd1 vccd1 vccd1 _3229_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5801_ _5798_/Y _5788_/Y _5799_/Y _5800_/X vssd1 vssd1 vccd1 vccd1 _5802_/A sky130_fd_sc_hd__o211ai_2
XFILLER_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5732_ _5556_/Y _5694_/X _5723_/Y _5731_/Y vssd1 vssd1 vccd1 vccd1 _5732_/Y sky130_fd_sc_hd__a2bb2oi_1
X_3993_ _3993_/A vssd1 vssd1 vccd1 vccd1 _4160_/C sky130_fd_sc_hd__clkbuf_2
X_5663_ _5663_/A _5663_/B _6002_/B _5842_/A vssd1 vssd1 vccd1 vccd1 _5825_/B sky130_fd_sc_hd__nand4_2
X_4614_ _4643_/A _4636_/A vssd1 vssd1 vccd1 vccd1 _4632_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5594_ _5594_/A _5842_/A vssd1 vssd1 vccd1 vccd1 _5604_/A sky130_fd_sc_hd__nand2_1
X_4545_ _4545_/A vssd1 vssd1 vccd1 vccd1 _4689_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4476_ _4476_/A _5534_/A _5678_/B vssd1 vssd1 vccd1 vccd1 _4476_/X sky130_fd_sc_hd__and3_1
X_6215_ _6222_/A _6214_/A _6214_/B vssd1 vssd1 vccd1 vccd1 _6215_/Y sky130_fd_sc_hd__o21ai_2
X_3427_ _3536_/A vssd1 vssd1 vccd1 vccd1 _3711_/A sky130_fd_sc_hd__clkbuf_2
X_6146_ _6164_/A _6180_/A _6164_/B vssd1 vssd1 vccd1 vccd1 _6148_/B sky130_fd_sc_hd__nand3_1
X_3358_ _3440_/A _4939_/A _5382_/C _3358_/D vssd1 vssd1 vccd1 vccd1 _3359_/C sky130_fd_sc_hd__nand4_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _6077_/A _6077_/B vssd1 vssd1 vccd1 vccd1 _6078_/B sky130_fd_sc_hd__nand2_1
X_3289_ _4026_/A vssd1 vssd1 vccd1 vccd1 _4540_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_45_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5028_ _4875_/A _4875_/B _4878_/A _4885_/A vssd1 vssd1 vccd1 vccd1 _5032_/B sky130_fd_sc_hd__a22oi_4
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4330_ _4333_/A _4330_/B vssd1 vssd1 vccd1 vccd1 _4331_/A sky130_fd_sc_hd__nand2_1
X_4261_ _4901_/B vssd1 vssd1 vccd1 vccd1 _4261_/Y sky130_fd_sc_hd__inv_2
X_3212_ _3458_/B _4366_/A vssd1 vssd1 vccd1 vccd1 _3215_/A sky130_fd_sc_hd__nand2_1
X_6000_ _6165_/B vssd1 vssd1 vccd1 vccd1 _6205_/C sky130_fd_sc_hd__clkbuf_2
X_4192_ _4936_/B vssd1 vssd1 vccd1 vccd1 _5925_/A sky130_fd_sc_hd__clkbuf_4
X_3143_ _3270_/B vssd1 vssd1 vccd1 vccd1 _3179_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3976_ _3976_/A _3976_/B _3976_/C vssd1 vssd1 vccd1 vccd1 _3977_/A sky130_fd_sc_hd__nand3_1
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5715_ _5719_/A _5933_/D _5719_/C _5719_/D vssd1 vssd1 vccd1 vccd1 _5729_/B sky130_fd_sc_hd__and4_1
XFILLER_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5646_ _5646_/A _5646_/B vssd1 vssd1 vccd1 vccd1 _5646_/Y sky130_fd_sc_hd__xnor2_2
X_5577_ _5404_/B _5918_/B _5919_/B _5580_/A vssd1 vssd1 vccd1 vccd1 _5654_/A sky130_fd_sc_hd__a22o_2
XFILLER_2_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4528_ _4532_/A _4935_/C vssd1 vssd1 vccd1 vccd1 _4529_/B sky130_fd_sc_hd__nand2_1
X_4459_ _4254_/B _4449_/Y _4458_/Y vssd1 vssd1 vccd1 vccd1 _4459_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6129_ _6132_/A _6132_/B _6236_/A _6235_/B vssd1 vssd1 vccd1 vccd1 _6129_/Y sky130_fd_sc_hd__o2bb2ai_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3830_ _3310_/B _3829_/C _6165_/A _4042_/B vssd1 vssd1 vccd1 vccd1 _3830_/Y sky130_fd_sc_hd__a22oi_4
X_3761_ _3761_/A _3761_/B vssd1 vssd1 vccd1 vccd1 _3761_/Y sky130_fd_sc_hd__nand2_1
X_5500_ _5497_/Y _5498_/X _5499_/Y vssd1 vssd1 vccd1 vccd1 _5514_/C sky130_fd_sc_hd__o21ai_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3692_ _4110_/B vssd1 vssd1 vccd1 vccd1 _5656_/A sky130_fd_sc_hd__buf_4
X_5431_ _5431_/A _5431_/B _5431_/C _5431_/D vssd1 vssd1 vccd1 vccd1 _5624_/A sky130_fd_sc_hd__nand4_2
X_5362_ _5184_/A _5184_/B _5184_/C _5195_/A _5520_/A vssd1 vssd1 vccd1 vccd1 _5363_/B
+ sky130_fd_sc_hd__a32oi_4
X_4313_ _4313_/A _4313_/B _4313_/C vssd1 vssd1 vccd1 vccd1 _4313_/X sky130_fd_sc_hd__and3_1
XFILLER_87_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5293_ _5128_/A _5120_/Y _5290_/Y _5292_/Y vssd1 vssd1 vccd1 vccd1 _5293_/Y sky130_fd_sc_hd__o2bb2ai_2
X_4244_ _4087_/Y _4088_/Y _4235_/Y _4236_/Y vssd1 vssd1 vccd1 vccd1 _4244_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4175_ _4137_/A _4137_/C _4137_/B _4141_/Y _4174_/Y vssd1 vssd1 vccd1 vccd1 _4315_/A
+ sky130_fd_sc_hd__a32oi_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3959_ _4935_/C vssd1 vssd1 vccd1 vccd1 _5792_/A sky130_fd_sc_hd__buf_4
X_5629_ _5629_/A _5634_/C _5634_/D vssd1 vssd1 vccd1 vccd1 _5631_/B sky130_fd_sc_hd__nand3_1
XFILLER_78_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5980_ _5980_/A _5980_/B _5980_/C vssd1 vssd1 vccd1 vccd1 _5981_/B sky130_fd_sc_hd__nand3_4
X_4931_ _4931_/A _5286_/A vssd1 vssd1 vccd1 vccd1 _4932_/B sky130_fd_sc_hd__nand2_2
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4862_ _5046_/A vssd1 vssd1 vccd1 vccd1 _5258_/A sky130_fd_sc_hd__buf_2
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3813_ _5511_/C _5858_/C _3814_/A vssd1 vssd1 vccd1 vccd1 _3813_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_15 _4849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4793_ _4801_/A _4801_/B _4796_/A _4796_/B vssd1 vssd1 vccd1 vccd1 _4793_/X sky130_fd_sc_hd__o2bb2a_2
X_3744_ _3603_/Y _3739_/Y _3743_/Y vssd1 vssd1 vccd1 vccd1 _3745_/B sky130_fd_sc_hd__o21ai_4
X_3675_ _4877_/A _3711_/A vssd1 vssd1 vccd1 vccd1 _3676_/B sky130_fd_sc_hd__nand2_2
X_5414_ _5263_/A _5249_/Y _5402_/Y _5405_/Y vssd1 vssd1 vccd1 vccd1 _5414_/Y sky130_fd_sc_hd__a22oi_4
X_5345_ _5340_/Y _5341_/Y _5342_/Y _5344_/Y vssd1 vssd1 vccd1 vccd1 _5364_/A sky130_fd_sc_hd__o211ai_4
X_5276_ _5272_/X _5273_/Y _5274_/Y _5275_/Y vssd1 vssd1 vccd1 vccd1 _5277_/C sky130_fd_sc_hd__o22ai_2
X_4227_ _4126_/Y _4127_/X _4130_/A _4130_/B vssd1 vssd1 vccd1 vccd1 _4227_/X sky130_fd_sc_hd__o22a_1
X_4158_ _3991_/A _3977_/A _4006_/Y vssd1 vssd1 vccd1 vccd1 _4159_/C sky130_fd_sc_hd__a21oi_1
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4089_ _4087_/Y _4088_/Y _4254_/A _3902_/B vssd1 vssd1 vccd1 vccd1 _4090_/A sky130_fd_sc_hd__o2bb2ai_1
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 a[7] vssd1 vssd1 vccd1 vccd1 _4906_/A sky130_fd_sc_hd__buf_2
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput24 b[17] vssd1 vssd1 vccd1 vccd1 _5230_/A sky130_fd_sc_hd__buf_4
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3460_ _3870_/A vssd1 vssd1 vccd1 vccd1 _4530_/A sky130_fd_sc_hd__clkbuf_4
X_3391_ _3483_/A _3382_/A _3483_/B vssd1 vssd1 vccd1 vccd1 _3392_/C sky130_fd_sc_hd__a21o_1
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5130_ _5130_/A _5130_/B _5130_/C vssd1 vssd1 vccd1 vccd1 _5131_/A sky130_fd_sc_hd__nand3_1
XFILLER_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5061_ _5081_/A _5081_/B _5060_/Y vssd1 vssd1 vccd1 vccd1 _5062_/C sky130_fd_sc_hd__a21o_1
X_4012_ _3985_/A _4009_/Y _3985_/B _4011_/X vssd1 vssd1 vccd1 vccd1 _4012_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_84_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5963_ _5960_/X _5961_/X _5962_/Y vssd1 vssd1 vccd1 vccd1 _5966_/A sky130_fd_sc_hd__o21ai_1
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4914_ _3634_/A _5453_/A _4776_/B _4907_/X _4903_/Y vssd1 vssd1 vccd1 vccd1 _4917_/B
+ sky130_fd_sc_hd__o221ai_4
X_5894_ _5892_/X _5893_/Y _5891_/A vssd1 vssd1 vccd1 vccd1 _5974_/D sky130_fd_sc_hd__o21bai_1
X_4845_ _4845_/A _4845_/B vssd1 vssd1 vccd1 vccd1 _5518_/A sky130_fd_sc_hd__nand2_2
X_4776_ _4776_/A _4776_/B vssd1 vssd1 vccd1 vccd1 _4784_/A sky130_fd_sc_hd__nand2_1
X_3727_ _6125_/A vssd1 vssd1 vccd1 vccd1 _3829_/C sky130_fd_sc_hd__buf_2
X_3658_ _3658_/A _3658_/B vssd1 vssd1 vccd1 vccd1 _3666_/B sky130_fd_sc_hd__nand2_1
X_3589_ _3593_/B _3593_/C _3592_/A vssd1 vssd1 vccd1 vccd1 _3591_/B sky130_fd_sc_hd__nand3_1
X_5328_ _5328_/A _5366_/C vssd1 vssd1 vccd1 vccd1 _5495_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5259_ _4860_/X _5603_/C _4868_/Y vssd1 vssd1 vccd1 vccd1 _5259_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4630_ _4630_/A _4630_/B _4635_/A _4635_/B vssd1 vssd1 vccd1 vccd1 _4631_/B sky130_fd_sc_hd__nand4_2
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4561_ _4367_/Y _4371_/Y _4377_/Y _4392_/Y vssd1 vssd1 vccd1 vccd1 _4561_/X sky130_fd_sc_hd__o211a_2
X_3512_ _5034_/A vssd1 vssd1 vccd1 vccd1 _3512_/X sky130_fd_sc_hd__buf_6
X_4492_ _4495_/A _4495_/B _4648_/A _4498_/C vssd1 vssd1 vccd1 vccd1 _4494_/B sky130_fd_sc_hd__nand4_2
X_6231_ _6233_/C vssd1 vssd1 vccd1 vccd1 _6255_/C sky130_fd_sc_hd__clkbuf_2
X_3443_ _4571_/B _4228_/A _4935_/B _4571_/A vssd1 vssd1 vccd1 vccd1 _3443_/X sky130_fd_sc_hd__a22o_2
X_6162_ _6118_/A _6118_/B _6219_/B vssd1 vssd1 vccd1 vccd1 _6163_/B sky130_fd_sc_hd__o21ai_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3215_/B _3342_/A _3345_/A _3354_/Y vssd1 vssd1 vccd1 vccd1 _3374_/X sky130_fd_sc_hd__o22a_1
X_5113_ _5113_/A _5113_/B vssd1 vssd1 vccd1 vccd1 _5113_/Y sky130_fd_sc_hd__nand2_1
X_6093_ _6094_/B _6149_/A _6094_/A vssd1 vssd1 vccd1 vccd1 _6097_/A sky130_fd_sc_hd__a21o_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5310_/A _5039_/Y _5043_/Y vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__a21oi_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5946_ _5940_/Y _5943_/Y _5944_/Y _5945_/Y vssd1 vssd1 vccd1 vccd1 _5948_/C sky130_fd_sc_hd__o2bb2ai_1
XFILLER_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5877_ _5912_/A vssd1 vssd1 vccd1 vccd1 _5877_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4828_ _5302_/B vssd1 vssd1 vccd1 vccd1 _4829_/A sky130_fd_sc_hd__buf_2
X_4759_ _4742_/X _4749_/Y _4757_/Y _4758_/X vssd1 vssd1 vccd1 vccd1 _4765_/A sky130_fd_sc_hd__o2bb2ai_1
XFILLER_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5800_ _5793_/Y _5794_/Y _5789_/Y vssd1 vssd1 vccd1 vccd1 _5800_/X sky130_fd_sc_hd__a21o_1
X_3992_ _4160_/A _4160_/B vssd1 vssd1 vccd1 vccd1 _3994_/A sky130_fd_sc_hd__nand2_1
X_5731_ _5725_/Y _5726_/Y _5727_/Y _5730_/Y vssd1 vssd1 vccd1 vccd1 _5731_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_22_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5662_ _5662_/A _5662_/B vssd1 vssd1 vccd1 vccd1 _5666_/A sky130_fd_sc_hd__nand2_1
X_4613_ _4609_/X _4610_/Y _4794_/A _4794_/B vssd1 vssd1 vccd1 vccd1 _4636_/A sky130_fd_sc_hd__o211ai_1
X_5593_ _5831_/B vssd1 vssd1 vccd1 vccd1 _6124_/B sky130_fd_sc_hd__clkbuf_2
X_4544_ _4832_/A _4541_/X _4543_/Y vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__a21oi_4
X_6214_ _6214_/A _6214_/B vssd1 vssd1 vccd1 vccd1 _6222_/B sky130_fd_sc_hd__or2_1
X_4475_ _5546_/A vssd1 vssd1 vccd1 vccd1 _5534_/A sky130_fd_sc_hd__clkbuf_4
X_3426_ _4430_/A vssd1 vssd1 vccd1 vccd1 _4571_/B sky130_fd_sc_hd__clkbuf_4
X_6145_ _6164_/A _6180_/A _6164_/B vssd1 vssd1 vccd1 vccd1 _6148_/A sky130_fd_sc_hd__a21o_1
X_3357_ _4184_/A vssd1 vssd1 vccd1 vccd1 _4939_/A sky130_fd_sc_hd__buf_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6076_/A _6076_/B vssd1 vssd1 vccd1 vccd1 _6078_/A sky130_fd_sc_hd__nand2_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5027_ _4779_/B _4080_/X _5025_/Y _5026_/Y vssd1 vssd1 vccd1 vccd1 _5032_/A sky130_fd_sc_hd__a22o_1
X_3288_ _3215_/B _3342_/A _5382_/C _4941_/A _3287_/X vssd1 vssd1 vccd1 vccd1 _3295_/B
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_38_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5929_ _5942_/C _5937_/A vssd1 vssd1 vccd1 vccd1 _5936_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4260_ _4260_/A vssd1 vssd1 vccd1 vccd1 _4901_/B sky130_fd_sc_hd__buf_2
X_3211_ _4026_/A vssd1 vssd1 vccd1 vccd1 _4366_/A sky130_fd_sc_hd__clkbuf_4
X_4191_ _4213_/A _4213_/B _4213_/C vssd1 vssd1 vccd1 vccd1 _4399_/A sky130_fd_sc_hd__and3_4
X_3142_ _3533_/B vssd1 vssd1 vccd1 vccd1 _3270_/B sky130_fd_sc_hd__buf_4
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3975_ _3975_/A _3975_/B vssd1 vssd1 vccd1 vccd1 _3976_/C sky130_fd_sc_hd__nand2_1
X_5714_ _5719_/C _5933_/D _5719_/D _5719_/A vssd1 vssd1 vccd1 vccd1 _5729_/A sky130_fd_sc_hd__a22oi_2
X_5645_ _5523_/A _5523_/B _5776_/A vssd1 vssd1 vccd1 vccd1 _5646_/B sky130_fd_sc_hd__o21ai_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5576_ _5662_/A vssd1 vssd1 vccd1 vccd1 _5674_/B sky130_fd_sc_hd__buf_2
X_4527_ _4502_/C _4502_/A _4526_/Y vssd1 vssd1 vccd1 vccd1 _4665_/A sky130_fd_sc_hd__a21o_1
X_4458_ _4593_/A _5285_/A vssd1 vssd1 vccd1 vccd1 _4458_/Y sky130_fd_sc_hd__nand2_1
X_3409_ _3366_/Y _3369_/Y _3362_/Y vssd1 vssd1 vccd1 vccd1 _3410_/B sky130_fd_sc_hd__a21oi_2
X_6128_ _6132_/A _6132_/B _6205_/C vssd1 vssd1 vccd1 vccd1 _6128_/Y sky130_fd_sc_hd__nand3_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4389_ _5134_/B vssd1 vssd1 vccd1 vccd1 _5302_/B sky130_fd_sc_hd__clkbuf_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6059_/A _6059_/B vssd1 vssd1 vccd1 vccd1 _6193_/B sky130_fd_sc_hd__nand2_2
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3760_ _4738_/A _4068_/A _4065_/A _4852_/A vssd1 vssd1 vccd1 vccd1 _3760_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5430_ _5430_/A _5614_/A _5614_/B _5614_/C vssd1 vssd1 vccd1 vccd1 _5431_/D sky130_fd_sc_hd__nand4_1
X_3691_ _3691_/A vssd1 vssd1 vccd1 vccd1 _3691_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5361_ _5520_/B _5517_/D vssd1 vssd1 vccd1 vccd1 _5363_/A sky130_fd_sc_hd__nand2_2
X_5292_ _5287_/A _5291_/X _5288_/Y vssd1 vssd1 vccd1 vccd1 _5292_/Y sky130_fd_sc_hd__o21ai_1
X_4312_ _4313_/B _4313_/C _4313_/A vssd1 vssd1 vccd1 vccd1 _4312_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4243_ _5132_/B _3620_/C _4236_/B _5399_/A _4230_/Y vssd1 vssd1 vccd1 vccd1 _4243_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4174_ _4174_/A _4174_/B vssd1 vssd1 vccd1 vccd1 _4174_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3958_ _5123_/B vssd1 vssd1 vccd1 vccd1 _4935_/C sky130_fd_sc_hd__clkbuf_2
X_3889_ _3889_/A vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__buf_2
X_5628_ _5628_/A vssd1 vssd1 vccd1 vccd1 _5634_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5559_ _5550_/Y _5556_/Y _5557_/Y _5558_/X vssd1 vssd1 vccd1 vccd1 _5567_/A sky130_fd_sc_hd__o211ai_4
XFILLER_4_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4930_ _4930_/A input2/X vssd1 vssd1 vccd1 vccd1 _5124_/A sky130_fd_sc_hd__nand2_4
XFILLER_17_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4861_ _4861_/A _5237_/A vssd1 vssd1 vccd1 vccd1 _5046_/A sky130_fd_sc_hd__nand2_1
X_3812_ _4422_/C vssd1 vssd1 vccd1 vccd1 _5511_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_16 _5197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4792_ _4792_/A vssd1 vssd1 vccd1 vccd1 _4796_/B sky130_fd_sc_hd__clkbuf_2
X_3743_ _6294_/A _3740_/Y _3853_/A _3998_/A _3742_/X vssd1 vssd1 vccd1 vccd1 _3743_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3674_ _3708_/A _3708_/B _3674_/C vssd1 vssd1 vccd1 vccd1 _3685_/B sky130_fd_sc_hd__nand3_2
X_5413_ _5413_/A _5413_/B _5413_/C vssd1 vssd1 vccd1 vccd1 _5614_/B sky130_fd_sc_hd__nand3_2
X_5344_ _5337_/X _5332_/B _5343_/X _5336_/Y vssd1 vssd1 vccd1 vccd1 _5344_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_87_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5275_ _5256_/B _5256_/C _5256_/A vssd1 vssd1 vccd1 vccd1 _5275_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4226_ _4313_/A _4226_/B _4313_/C vssd1 vssd1 vccd1 vccd1 _4321_/B sky130_fd_sc_hd__nand3_2
X_4157_ _4157_/A _4157_/B _4157_/C vssd1 vssd1 vccd1 vccd1 _4159_/B sky130_fd_sc_hd__nand3_1
X_4088_ _4877_/A _4234_/A vssd1 vssd1 vccd1 vccd1 _4088_/Y sky130_fd_sc_hd__nand2_2
XFILLER_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput25 b[18] vssd1 vssd1 vccd1 vccd1 _5238_/A sky130_fd_sc_hd__clkbuf_4
Xinput14 a[8] vssd1 vssd1 vccd1 vccd1 _3510_/A sky130_fd_sc_hd__clkbuf_4
X_3390_ _3484_/A _3483_/B _3483_/A vssd1 vssd1 vccd1 vccd1 _3392_/B sky130_fd_sc_hd__nand3_1
X_5060_ _5229_/A _5658_/A vssd1 vssd1 vccd1 vccd1 _5060_/Y sky130_fd_sc_hd__nand2_2
X_4011_ _4157_/C _4011_/B vssd1 vssd1 vccd1 vccd1 _4011_/X sky130_fd_sc_hd__and2b_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5962_ _5865_/C _5865_/B _5829_/X vssd1 vssd1 vccd1 vccd1 _5962_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4913_ _4917_/A _4913_/B _4913_/C vssd1 vssd1 vccd1 vccd1 _4922_/A sky130_fd_sc_hd__nand3b_1
X_5893_ _5892_/B _5892_/C _5892_/A vssd1 vssd1 vccd1 vccd1 _5893_/Y sky130_fd_sc_hd__a21oi_1
X_4844_ _4845_/A _4845_/B _5980_/A vssd1 vssd1 vccd1 vccd1 _4848_/A sky130_fd_sc_hd__a21o_1
XFILLER_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4775_ _5207_/A _5286_/B vssd1 vssd1 vccd1 vccd1 _4776_/B sky130_fd_sc_hd__nand2_2
X_3726_ _5794_/A vssd1 vssd1 vccd1 vccd1 _6125_/A sky130_fd_sc_hd__buf_2
X_3657_ _3657_/A _3657_/B vssd1 vssd1 vccd1 vccd1 _3658_/B sky130_fd_sc_hd__nand2_1
X_3588_ _3482_/A _3593_/C _3592_/A vssd1 vssd1 vccd1 vccd1 _3591_/A sky130_fd_sc_hd__a21o_1
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5327_ _5366_/D vssd1 vssd1 vccd1 vccd1 _5327_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5258_ _5258_/A vssd1 vssd1 vccd1 vccd1 _5603_/C sky130_fd_sc_hd__clkbuf_4
X_5189_ _5189_/A _5189_/B _5189_/C vssd1 vssd1 vccd1 vccd1 _5520_/A sky130_fd_sc_hd__nand3_4
XFILLER_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4209_ _4516_/C _4209_/B vssd1 vssd1 vccd1 vccd1 _4219_/B sky130_fd_sc_hd__nor2_1
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4560_ _4560_/A vssd1 vssd1 vccd1 vccd1 _4817_/A sky130_fd_sc_hd__clkbuf_2
X_4491_ _4647_/B vssd1 vssd1 vccd1 vccd1 _4498_/C sky130_fd_sc_hd__clkbuf_2
X_3511_ _3633_/A vssd1 vssd1 vccd1 vccd1 _5034_/A sky130_fd_sc_hd__clkbuf_4
X_6230_ _6230_/A vssd1 vssd1 vccd1 vccd1 _6247_/B sky130_fd_sc_hd__inv_2
X_3442_ _3870_/A vssd1 vssd1 vccd1 vccd1 _3448_/A sky130_fd_sc_hd__inv_2
X_6161_ _6161_/A _6161_/B vssd1 vssd1 vccd1 vccd1 _6219_/A sky130_fd_sc_hd__nor2_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _3306_/Y _3300_/C _3305_/Y _3304_/Y vssd1 vssd1 vccd1 vccd1 _3398_/B sky130_fd_sc_hd__o2bb2ai_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5278_/A _5202_/B _5203_/A vssd1 vssd1 vccd1 vccd1 _5116_/B sky130_fd_sc_hd__nand3_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6091_/Y _6023_/C _6091_/B vssd1 vssd1 vccd1 vccd1 _6094_/A sky130_fd_sc_hd__o21ai_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5310_/A _5309_/A _5309_/B vssd1 vssd1 vccd1 vccd1 _5043_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_84_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5945_ _5945_/A vssd1 vssd1 vccd1 vccd1 _5945_/Y sky130_fd_sc_hd__inv_2
X_5876_ _5829_/X _5957_/B _5863_/X _5870_/Y vssd1 vssd1 vccd1 vccd1 _5879_/B sky130_fd_sc_hd__o211ai_1
X_4827_ _4827_/A _5006_/A _5506_/A _5348_/D vssd1 vssd1 vccd1 vccd1 _4827_/X sky130_fd_sc_hd__and4_1
X_4758_ _4890_/A _4890_/B _4758_/C vssd1 vssd1 vccd1 vccd1 _4758_/X sky130_fd_sc_hd__and3_1
X_3709_ _3684_/A _3684_/B _3707_/X _3708_/Y _3667_/X vssd1 vssd1 vccd1 vccd1 _3719_/B
+ sky130_fd_sc_hd__o221ai_2
X_4689_ _4689_/A _4689_/B vssd1 vssd1 vccd1 vccd1 _4689_/X sky130_fd_sc_hd__and2_1
XFILLER_0_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3991_ _3991_/A _4160_/A _4160_/B vssd1 vssd1 vccd1 vccd1 _3996_/C sky130_fd_sc_hd__nand3_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5730_ _5730_/A _5730_/B vssd1 vssd1 vccd1 vccd1 _5730_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5661_ _5661_/A _5661_/B vssd1 vssd1 vccd1 vccd1 _5661_/Y sky130_fd_sc_hd__nand2_1
X_4612_ _4606_/B _4606_/C _4599_/B vssd1 vssd1 vccd1 vccd1 _4794_/B sky130_fd_sc_hd__a21o_1
X_5592_ _5678_/A _5676_/A _5681_/A _5596_/A vssd1 vssd1 vccd1 vccd1 _5592_/Y sky130_fd_sc_hd__a22oi_2
X_4543_ _4539_/A _4540_/Y _4542_/Y vssd1 vssd1 vccd1 vccd1 _4543_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6213_ _6213_/A _6228_/A vssd1 vssd1 vccd1 vccd1 _6214_/B sky130_fd_sc_hd__xnor2_1
X_4474_ _4257_/Y _4473_/X _4459_/Y vssd1 vssd1 vccd1 vccd1 _4474_/Y sky130_fd_sc_hd__a21oi_1
X_3425_ input7/X vssd1 vssd1 vccd1 vccd1 _4430_/A sky130_fd_sc_hd__buf_2
X_6144_ _6089_/A _6089_/C _6089_/B vssd1 vssd1 vccd1 vccd1 _6164_/B sky130_fd_sc_hd__a21bo_1
XFILLER_38_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3356_ _3356_/A vssd1 vssd1 vccd1 vccd1 _4184_/A sky130_fd_sc_hd__clkbuf_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6170_/A _6076_/A _6076_/B _6077_/B vssd1 vssd1 vccd1 vccd1 _6081_/A sky130_fd_sc_hd__nand4_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3287_ _3287_/A vssd1 vssd1 vccd1 vccd1 _3287_/X sky130_fd_sc_hd__clkbuf_2
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5026_/A _5026_/B _5212_/B _5539_/B vssd1 vssd1 vccd1 vccd1 _5026_/Y sky130_fd_sc_hd__nand4_4
XFILLER_65_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5928_ _5926_/Y _5927_/X _6025_/C vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__o21bai_2
X_5859_ _5860_/B _5860_/C _5672_/X _5685_/X vssd1 vssd1 vccd1 vccd1 _5859_/Y sky130_fd_sc_hd__o2bb2ai_2
XFILLER_21_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3210_ _3210_/A vssd1 vssd1 vccd1 vccd1 _4026_/A sky130_fd_sc_hd__clkbuf_2
X_4190_ _4186_/Y _4189_/Y _4023_/Y vssd1 vssd1 vccd1 vccd1 _4213_/C sky130_fd_sc_hd__o21ai_1
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3141_ input7/X vssd1 vssd1 vccd1 vccd1 _3533_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_94_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3974_ _4152_/A _4011_/B vssd1 vssd1 vccd1 vccd1 _3975_/B sky130_fd_sc_hd__nand2_1
X_5713_ _5808_/A _5808_/B _5986_/B _5534_/A vssd1 vssd1 vccd1 vccd1 _5719_/A sky130_fd_sc_hd__a22o_1
X_5644_ _5776_/C _5776_/D vssd1 vssd1 vccd1 vccd1 _5646_/A sky130_fd_sc_hd__nand2_1
X_5575_ _5575_/A _5575_/B vssd1 vssd1 vccd1 vccd1 _5662_/A sky130_fd_sc_hd__nand2_2
X_4526_ _4494_/B _4494_/C _4494_/A vssd1 vssd1 vccd1 vccd1 _4526_/Y sky130_fd_sc_hd__a21oi_2
X_4457_ _4463_/A _4463_/B _4451_/X _4456_/X vssd1 vssd1 vccd1 vccd1 _4466_/A sky130_fd_sc_hd__o2bb2ai_2
X_3408_ _3402_/Y _3498_/A _3407_/X vssd1 vssd1 vccd1 vccd1 _3410_/A sky130_fd_sc_hd__o21ai_2
XFILLER_85_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4388_ _3186_/A _4711_/C _4362_/B vssd1 vssd1 vccd1 vccd1 _4680_/B sky130_fd_sc_hd__o21ai_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ _6127_/A _6127_/B _6127_/C _6127_/D vssd1 vssd1 vccd1 vccd1 _6132_/B sky130_fd_sc_hd__nand4_4
X_3339_ _3533_/A _5053_/A _4369_/A _3542_/A vssd1 vssd1 vccd1 vccd1 _3348_/B sky130_fd_sc_hd__nand4_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _6058_/A _6058_/B _6058_/C _6058_/D vssd1 vssd1 vccd1 vccd1 _6059_/B sky130_fd_sc_hd__nand4_1
XFILLER_73_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5009_ _5001_/Y _5005_/Y _5008_/Y _4711_/D vssd1 vssd1 vccd1 vccd1 _5012_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_26_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3690_ _3699_/A _3699_/B _3689_/A vssd1 vssd1 vccd1 vccd1 _3690_/Y sky130_fd_sc_hd__a21oi_2
X_5360_ _5519_/A _5519_/B _5519_/C vssd1 vssd1 vccd1 vccd1 _5517_/D sky130_fd_sc_hd__nand3_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5291_ _5291_/A vssd1 vssd1 vccd1 vccd1 _5291_/X sky130_fd_sc_hd__clkbuf_2
X_4311_ _4313_/A _4224_/X _4321_/B _4322_/B _4322_/A vssd1 vssd1 vccd1 vccd1 _4315_/B
+ sky130_fd_sc_hd__o2111ai_2
X_4242_ _4231_/Y _4232_/Y _4237_/X _4241_/X vssd1 vssd1 vccd1 vccd1 _4302_/C sky130_fd_sc_hd__o211ai_4
XFILLER_95_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4173_ _3968_/A _4143_/X _4054_/A _4054_/B vssd1 vssd1 vccd1 vccd1 _4174_/B sky130_fd_sc_hd__o211ai_1
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3957_ _3803_/A _5919_/A _5442_/C _4201_/A vssd1 vssd1 vccd1 vccd1 _3964_/A sky130_fd_sc_hd__a22o_1
X_3888_ _4430_/A _4906_/B vssd1 vssd1 vccd1 vccd1 _3889_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5627_ _5627_/A _5627_/B _5627_/C vssd1 vssd1 vccd1 vccd1 _5628_/A sky130_fd_sc_hd__nand3_1
X_5558_ _5561_/C _5694_/C _5550_/A vssd1 vssd1 vccd1 vccd1 _5558_/X sky130_fd_sc_hd__a21o_1
X_4509_ _4502_/A _4502_/B _4502_/C vssd1 vssd1 vccd1 vccd1 _4511_/A sky130_fd_sc_hd__a21oi_1
X_5489_ _5489_/A _5614_/B _5614_/C vssd1 vssd1 vccd1 vccd1 _5490_/C sky130_fd_sc_hd__nand3_1
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _4860_/A vssd1 vssd1 vccd1 vccd1 _4860_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3811_ _3667_/X _3685_/C _3685_/B vssd1 vssd1 vccd1 vccd1 _3811_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4791_ _4950_/A _4951_/A _4950_/B vssd1 vssd1 vccd1 vccd1 _4792_/A sky130_fd_sc_hd__and3_1
XANTENNA_17 _5230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3742_ _3609_/X _3610_/Y _3733_/Y _3734_/X vssd1 vssd1 vccd1 vccd1 _3742_/X sky130_fd_sc_hd__a2bb2o_1
X_3673_ _3530_/B _3747_/A _5382_/C _4621_/C _3761_/A vssd1 vssd1 vccd1 vccd1 _3674_/C
+ sky130_fd_sc_hd__o2111ai_2
X_5412_ _5208_/Y _5212_/X _5411_/X vssd1 vssd1 vccd1 vccd1 _5413_/C sky130_fd_sc_hd__a21oi_4
X_5343_ _5143_/Y _5139_/Y _5142_/X _5152_/X _4965_/X vssd1 vssd1 vccd1 vccd1 _5343_/X
+ sky130_fd_sc_hd__o32a_1
X_5274_ _5424_/A _5424_/B _5269_/A vssd1 vssd1 vccd1 vccd1 _5274_/Y sky130_fd_sc_hd__a21oi_1
X_4225_ _4225_/A vssd1 vssd1 vccd1 vccd1 _4313_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4156_ _4157_/A _4151_/A _4157_/C vssd1 vssd1 vccd1 vccd1 _4159_/A sky130_fd_sc_hd__a21o_1
XFILLER_28_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4087_ _5065_/A _4931_/A vssd1 vssd1 vccd1 vccd1 _4087_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4989_ _4989_/A _4989_/B vssd1 vssd1 vccd1 vccd1 _4989_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput15 a[9] vssd1 vssd1 vccd1 vccd1 _3952_/A sky130_fd_sc_hd__clkbuf_2
Xinput26 b[1] vssd1 vssd1 vccd1 vccd1 _3473_/A sky130_fd_sc_hd__buf_4
X_4010_ _4010_/A _4052_/A _4010_/C vssd1 vssd1 vccd1 vccd1 _4157_/C sky130_fd_sc_hd__nor3_2
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5961_ _5877_/X _5869_/Y _5900_/Y _5956_/B vssd1 vssd1 vccd1 vccd1 _5961_/X sky130_fd_sc_hd__o211a_1
XFILLER_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4912_ _4909_/Y _4917_/A _4918_/A vssd1 vssd1 vccd1 vccd1 _4912_/Y sky130_fd_sc_hd__a21boi_2
X_5892_ _5892_/A _5892_/B _5892_/C vssd1 vssd1 vccd1 vccd1 _5892_/X sky130_fd_sc_hd__and3_1
XFILLER_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4843_ _4840_/X _4841_/X _4842_/Y _4523_/S vssd1 vssd1 vccd1 vccd1 _5980_/A sky130_fd_sc_hd__o22ai_4
XFILLER_33_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4774_ _5026_/B _4777_/C vssd1 vssd1 vccd1 vccd1 _4776_/A sky130_fd_sc_hd__nand2_1
X_3725_ _5286_/A vssd1 vssd1 vccd1 vccd1 _5794_/A sky130_fd_sc_hd__clkbuf_4
X_3656_ _3656_/A _3707_/C vssd1 vssd1 vccd1 vccd1 _3666_/A sky130_fd_sc_hd__nand2_1
X_3587_ _3857_/A _3853_/A vssd1 vssd1 vccd1 vccd1 _3601_/A sky130_fd_sc_hd__nand2_1
X_5326_ _5277_/Y _5283_/Y _5320_/Y _5321_/X vssd1 vssd1 vccd1 vccd1 _5331_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5257_ _5257_/A _5257_/B vssd1 vssd1 vccd1 vccd1 _5257_/Y sky130_fd_sc_hd__nand2_1
X_4208_ _3639_/B _6077_/A _6076_/B _4362_/C vssd1 vssd1 vccd1 vccd1 _4209_/B sky130_fd_sc_hd__a22oi_4
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5188_ _5019_/Y _5005_/Y _5020_/Y _5021_/X vssd1 vssd1 vccd1 vccd1 _5189_/C sky130_fd_sc_hd__o2bb2ai_1
X_4139_ _4134_/Y _4135_/X _4130_/Y _4131_/Y vssd1 vssd1 vccd1 vccd1 _4141_/B sky130_fd_sc_hd__o22ai_2
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3510_ _3510_/A vssd1 vssd1 vccd1 vccd1 _3633_/A sky130_fd_sc_hd__inv_2
X_4490_ _4490_/A _4490_/B _4490_/C vssd1 vssd1 vccd1 vccd1 _4647_/B sky130_fd_sc_hd__nand3_1
X_3441_ _3441_/A vssd1 vssd1 vccd1 vccd1 _3441_/X sky130_fd_sc_hd__buf_4
X_6160_ _6110_/D _6159_/Y _6156_/Y _6157_/X vssd1 vssd1 vccd1 vccd1 _6161_/B sky130_fd_sc_hd__a22oi_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3372_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3398_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5111_ _5278_/A _5203_/A _5202_/B vssd1 vssd1 vccd1 vccd1 _5116_/A sky130_fd_sc_hd__a21o_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6091_/A _6091_/B vssd1 vssd1 vccd1 vccd1 _6091_/Y sky130_fd_sc_hd__nand2_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5042_/A vssd1 vssd1 vccd1 vccd1 _5309_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5944_ _5944_/A _5944_/B vssd1 vssd1 vccd1 vccd1 _5944_/Y sky130_fd_sc_hd__nor2_1
X_5875_ _5786_/B _5873_/X _5874_/Y vssd1 vssd1 vccd1 vccd1 _5879_/A sky130_fd_sc_hd__o21ai_1
X_4826_ _6233_/A vssd1 vssd1 vccd1 vccd1 _5506_/A sky130_fd_sc_hd__buf_2
XFILLER_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4757_ _4890_/A _4890_/B _4758_/C vssd1 vssd1 vccd1 vccd1 _4757_/Y sky130_fd_sc_hd__a21oi_2
X_4688_ _4661_/A _4661_/B _4661_/C _4663_/A _4669_/Y vssd1 vssd1 vccd1 vccd1 _4819_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3708_ _3708_/A _3708_/B vssd1 vssd1 vccd1 vccd1 _3708_/Y sky130_fd_sc_hd__nand2_1
X_3639_ _3639_/A _3639_/B _5850_/A _5905_/B vssd1 vssd1 vccd1 vccd1 _3639_/X sky130_fd_sc_hd__and4_2
X_5309_ _5309_/A _5309_/B vssd1 vssd1 vccd1 vccd1 _5310_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6289_ _6289_/A _6289_/B _6289_/C vssd1 vssd1 vccd1 vccd1 _6290_/B sky130_fd_sc_hd__and3_1
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3990_ _3990_/A _3990_/B _3990_/C vssd1 vssd1 vccd1 vccd1 _4160_/B sky130_fd_sc_hd__nand3_2
XFILLER_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5660_ _5598_/A _5598_/B _5604_/A vssd1 vssd1 vccd1 vccd1 _5661_/B sky130_fd_sc_hd__o21ai_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4611_ _4574_/Y _4577_/Y _4606_/C _4599_/B vssd1 vssd1 vccd1 vccd1 _4794_/A sky130_fd_sc_hd__o211ai_1
X_5591_ _5608_/A _5608_/B _5608_/C vssd1 vssd1 vccd1 vccd1 _5686_/A sky130_fd_sc_hd__nand3_1
X_4542_ _4542_/A _5302_/B vssd1 vssd1 vccd1 vccd1 _4542_/Y sky130_fd_sc_hd__nand2_1
X_4473_ _4592_/A vssd1 vssd1 vccd1 vccd1 _4473_/X sky130_fd_sc_hd__clkbuf_2
X_6212_ _6212_/A _6212_/B vssd1 vssd1 vccd1 vccd1 _6228_/A sky130_fd_sc_hd__nor2_1
X_3424_ _3419_/Y _3421_/Y _3423_/Y vssd1 vssd1 vccd1 vccd1 _3465_/B sky130_fd_sc_hd__a21o_1
X_6143_ _6143_/A _6143_/B _6143_/C vssd1 vssd1 vccd1 vccd1 _6180_/A sky130_fd_sc_hd__nand3_2
X_3355_ _3345_/A _3354_/Y _3345_/B vssd1 vssd1 vccd1 vccd1 _3359_/B sky130_fd_sc_hd__o21ai_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _5240_/B vssd1 vssd1 vccd1 vccd1 _5382_/C sky130_fd_sc_hd__clkbuf_4
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6236_/A _6072_/Y _6073_/X _6069_/Y vssd1 vssd1 vccd1 vccd1 _6089_/B sky130_fd_sc_hd__o211ai_4
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5025_/A _5025_/B vssd1 vssd1 vccd1 vccd1 _5025_/Y sky130_fd_sc_hd__nand2_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5927_ _5927_/A _5927_/B _5927_/C vssd1 vssd1 vccd1 vccd1 _5927_/X sky130_fd_sc_hd__and3_1
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5858_ _5868_/A _5868_/B _5858_/C _6205_/B vssd1 vssd1 vccd1 vccd1 _5860_/C sky130_fd_sc_hd__nand4_4
X_5789_ _5925_/A _5931_/A vssd1 vssd1 vccd1 vccd1 _5789_/Y sky130_fd_sc_hd__nand2_1
X_4809_ _4809_/A _4809_/B vssd1 vssd1 vccd1 vccd1 _4814_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3140_ _3140_/A vssd1 vssd1 vccd1 vccd1 _3150_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_79_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5712_ _5712_/A _5933_/C _6016_/A _5986_/B vssd1 vssd1 vccd1 vccd1 _5719_/D sky130_fd_sc_hd__nand4_2
X_3973_ _3973_/A _3973_/B vssd1 vssd1 vccd1 vccd1 _3975_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5643_ _5643_/A _5643_/B _5643_/C _5643_/D vssd1 vssd1 vccd1 vccd1 _5776_/D sky130_fd_sc_hd__nand4_1
X_5574_ _5246_/X _5598_/A _5571_/Y _5573_/Y vssd1 vssd1 vccd1 vccd1 _5584_/A sky130_fd_sc_hd__o22a_2
X_4525_ _4681_/A _4681_/B _4516_/B vssd1 vssd1 vccd1 vccd1 _4525_/X sky130_fd_sc_hd__o21a_1
X_4456_ _4453_/Y _4456_/B _4890_/C _5546_/A vssd1 vssd1 vccd1 vccd1 _4456_/X sky130_fd_sc_hd__and4b_1
XFILLER_49_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3407_ _4542_/A _5663_/A _5663_/B _4390_/A vssd1 vssd1 vccd1 vccd1 _3407_/X sky130_fd_sc_hd__a22o_1
X_4387_ _4387_/A vssd1 vssd1 vccd1 vccd1 _4711_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_58_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3338_ _3536_/A vssd1 vssd1 vccd1 vccd1 _3542_/A sky130_fd_sc_hd__buf_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6126_ _6236_/C _6126_/B vssd1 vssd1 vccd1 vccd1 _6132_/A sky130_fd_sc_hd__nand2_1
XFILLER_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _5966_/A _5966_/B _5966_/C _5969_/C vssd1 vssd1 vccd1 vccd1 _6058_/D sky130_fd_sc_hd__a31o_1
X_3269_ _3870_/A vssd1 vssd1 vccd1 vccd1 _4958_/B sky130_fd_sc_hd__buf_4
X_5008_ _5006_/Y _5007_/Y _4711_/A _4674_/X vssd1 vssd1 vccd1 vccd1 _5008_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_45_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5290_ _5794_/A _4080_/X _5794_/B _5546_/A vssd1 vssd1 vccd1 vccd1 _5290_/Y sky130_fd_sc_hd__a22oi_4
X_4310_ _4310_/A vssd1 vssd1 vccd1 vccd1 _4322_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4241_ _4238_/Y _4422_/A _4230_/Y vssd1 vssd1 vccd1 vccd1 _4241_/X sky130_fd_sc_hd__a21o_2
XFILLER_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4172_ _4054_/A _4054_/B _4054_/C vssd1 vssd1 vccd1 vccd1 _4174_/A sky130_fd_sc_hd__a21bo_1
XFILLER_67_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3956_ _5284_/D vssd1 vssd1 vccd1 vccd1 _5442_/C sky130_fd_sc_hd__buf_4
X_5626_ _5566_/A _5568_/A _5625_/C _5625_/D vssd1 vssd1 vccd1 vccd1 _5627_/C sky130_fd_sc_hd__a22o_1
X_3887_ _4260_/A vssd1 vssd1 vccd1 vccd1 _4906_/B sky130_fd_sc_hd__clkbuf_2
X_5557_ _5413_/B _5413_/C _5414_/Y vssd1 vssd1 vccd1 vccd1 _5557_/Y sky130_fd_sc_hd__a21oi_2
X_5488_ _5484_/Y _5485_/Y _5486_/Y _5487_/Y vssd1 vssd1 vccd1 vccd1 _5493_/A sky130_fd_sc_hd__o22ai_1
X_4508_ _4506_/C _4506_/B _4506_/A vssd1 vssd1 vccd1 vccd1 _4508_/Y sky130_fd_sc_hd__a21oi_2
X_4439_ _5539_/B vssd1 vssd1 vccd1 vccd1 _5931_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6109_ _6110_/A _6110_/B _6159_/A _6110_/D vssd1 vssd1 vccd1 vccd1 _6112_/A sky130_fd_sc_hd__a22o_1
XFILLER_58_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3810_ _3810_/A _3810_/B vssd1 vssd1 vccd1 vccd1 _3810_/Y sky130_fd_sc_hd__nor2_2
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4790_ _4950_/A _4951_/A _4950_/B vssd1 vssd1 vccd1 vccd1 _4796_/A sky130_fd_sc_hd__a21oi_4
X_3741_ _3736_/X _3737_/Y _3733_/Y _3734_/X vssd1 vssd1 vccd1 vccd1 _3998_/A sky130_fd_sc_hd__o211ai_4
XANTENNA_18 _5230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3672_ _5299_/B vssd1 vssd1 vccd1 vccd1 _4621_/C sky130_fd_sc_hd__buf_4
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5411_ _5833_/A _5663_/B _5411_/C _5688_/A vssd1 vssd1 vccd1 vccd1 _5411_/X sky130_fd_sc_hd__and4_4
X_5342_ _5170_/B _5171_/C _5177_/Y _5178_/Y vssd1 vssd1 vccd1 vccd1 _5342_/Y sky130_fd_sc_hd__o2bb2ai_2
X_5273_ _5224_/Y _5026_/Y _5281_/A _5281_/B _5220_/Y vssd1 vssd1 vccd1 vccd1 _5273_/Y
+ sky130_fd_sc_hd__a221oi_2
X_4224_ _4313_/B _4225_/A _4224_/C vssd1 vssd1 vccd1 vccd1 _4224_/X sky130_fd_sc_hd__and3_1
X_4155_ _4006_/Y _4007_/Y _4152_/Y _4154_/Y vssd1 vssd1 vccd1 vccd1 _4166_/B sky130_fd_sc_hd__o211ai_4
XFILLER_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4086_ _3474_/A _3669_/X _3902_/B _4254_/A _4085_/X vssd1 vssd1 vccd1 vccd1 _4091_/A
+ sky130_fd_sc_hd__o221ai_4
XFILLER_36_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4988_ _4988_/A _4988_/B _4988_/C _4988_/D vssd1 vssd1 vccd1 vccd1 _4989_/B sky130_fd_sc_hd__nand4_1
X_3939_ _3939_/A _3946_/A vssd1 vssd1 vccd1 vccd1 _3985_/B sky130_fd_sc_hd__nand2_1
X_5609_ _5686_/B _5609_/B vssd1 vssd1 vccd1 vccd1 _5609_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 b[0] vssd1 vssd1 vccd1 vccd1 _4176_/A sky130_fd_sc_hd__buf_4
Xinput27 b[2] vssd1 vssd1 vccd1 vccd1 _3256_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5960_ _5960_/A _5960_/B _5960_/C vssd1 vssd1 vccd1 vccd1 _5960_/X sky130_fd_sc_hd__and3_1
XFILLER_80_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5891_ _5891_/A _5891_/B _5891_/C vssd1 vssd1 vccd1 vccd1 _5974_/C sky130_fd_sc_hd__nand3_1
X_4911_ _4779_/Y _4784_/B _4784_/A vssd1 vssd1 vccd1 vccd1 _4918_/A sky130_fd_sc_hd__a21boi_2
XFILLER_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4842_ _4842_/A _4842_/B _4842_/C _4842_/D vssd1 vssd1 vccd1 vccd1 _4842_/Y sky130_fd_sc_hd__nand4_2
XFILLER_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4773_ _4473_/X _4592_/B _4593_/Y _4589_/Y vssd1 vssd1 vccd1 vccd1 _4781_/A sky130_fd_sc_hd__o22a_1
X_3724_ _3952_/A vssd1 vssd1 vccd1 vccd1 _5286_/A sky130_fd_sc_hd__buf_2
X_3655_ _5229_/A _4423_/A vssd1 vssd1 vccd1 vccd1 _3707_/C sky130_fd_sc_hd__and2_1
X_3586_ _3586_/A _3586_/B _3586_/C vssd1 vssd1 vccd1 vccd1 _3853_/A sky130_fd_sc_hd__nand3_2
X_5325_ _5325_/A _5325_/B vssd1 vssd1 vccd1 vccd1 _5331_/A sky130_fd_sc_hd__nand2_1
X_5256_ _5256_/A _5256_/B _5256_/C vssd1 vssd1 vccd1 vccd1 _5490_/A sky130_fd_sc_hd__nand3_2
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4207_ _5809_/B vssd1 vssd1 vccd1 vccd1 _6076_/B sky130_fd_sc_hd__clkbuf_4
X_5187_ _4956_/X _4958_/X _4943_/C _5182_/A _5182_/B vssd1 vssd1 vccd1 vccd1 _5189_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_68_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4138_ _4053_/Y _4054_/X _4123_/Y _4125_/Y _4317_/A vssd1 vssd1 vccd1 vccd1 _4138_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4069_ _5240_/B _5285_/A vssd1 vssd1 vccd1 vccd1 _4069_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3440_ _3440_/A _3440_/B vssd1 vssd1 vccd1 vccd1 _3445_/B sky130_fd_sc_hd__nand2_1
X_3371_ _3362_/Y _3367_/Y _3370_/X vssd1 vssd1 vccd1 vccd1 _3372_/B sky130_fd_sc_hd__o21ai_2
X_6090_ _6090_/A _6090_/B _6090_/C vssd1 vssd1 vccd1 vccd1 _6149_/A sky130_fd_sc_hd__nand3_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5110_/A _5110_/B vssd1 vssd1 vccd1 vccd1 _5202_/B sky130_fd_sc_hd__nand2_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5041_ _5032_/B _5041_/B _5041_/C vssd1 vssd1 vccd1 vccd1 _5309_/A sky130_fd_sc_hd__nand3b_2
XFILLER_84_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5943_ _5940_/C _5943_/B _5943_/C vssd1 vssd1 vccd1 vccd1 _5943_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5874_ _5860_/A _5786_/Y _5732_/Y _5740_/X vssd1 vssd1 vccd1 vccd1 _5874_/Y sky130_fd_sc_hd__o22ai_1
X_4825_ _4832_/A _4687_/Y _4819_/Y _4824_/Y vssd1 vssd1 vccd1 vccd1 _5190_/A sky130_fd_sc_hd__a22oi_1
XFILLER_21_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4756_ _5064_/A _5448_/B vssd1 vssd1 vccd1 vccd1 _4758_/C sky130_fd_sc_hd__and2_1
X_3707_ _3761_/A _3754_/B _3707_/C vssd1 vssd1 vccd1 vccd1 _3707_/X sky130_fd_sc_hd__and3_1
X_4687_ _3473_/Y _4674_/X _4540_/Y vssd1 vssd1 vccd1 vccd1 _4687_/Y sky130_fd_sc_hd__o21ai_1
X_3638_ _5663_/B vssd1 vssd1 vccd1 vccd1 _5905_/B sky130_fd_sc_hd__clkbuf_2
X_3569_ _3576_/A _3730_/B _3577_/B _3703_/B vssd1 vssd1 vccd1 vccd1 _3736_/A sky130_fd_sc_hd__a22o_1
X_5308_ _5321_/B vssd1 vssd1 vccd1 vccd1 _5366_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6288_ _6289_/B _6289_/C _6289_/A vssd1 vssd1 vccd1 vccd1 _6290_/A sky130_fd_sc_hd__a21oi_1
XFILLER_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5239_ _4277_/C _5831_/B _5677_/A _3270_/B vssd1 vssd1 vccd1 vccd1 _5239_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4610_ _4601_/B _4441_/C _4601_/A _4463_/C vssd1 vssd1 vccd1 vccd1 _4610_/Y sky130_fd_sc_hd__a31oi_1
X_5590_ _5608_/B _5608_/C _5608_/A vssd1 vssd1 vccd1 vccd1 _5590_/Y sky130_fd_sc_hd__a21oi_2
X_4541_ _3473_/Y _4387_/A _4540_/Y vssd1 vssd1 vccd1 vccd1 _4541_/X sky130_fd_sc_hd__o21a_1
X_4472_ _4453_/Y _4459_/Y _4461_/Y _4463_/B _4463_/A vssd1 vssd1 vccd1 vccd1 _4640_/A
+ sky130_fd_sc_hd__o2111ai_4
X_6211_ _6240_/D _6240_/C _6240_/B _6227_/A _6183_/A vssd1 vssd1 vccd1 vccd1 _6212_/B
+ sky130_fd_sc_hd__a311oi_1
X_3423_ _4193_/A _4236_/A vssd1 vssd1 vccd1 vccd1 _3423_/Y sky130_fd_sc_hd__nand2_1
X_6142_ _6143_/A _6143_/B _6143_/C vssd1 vssd1 vccd1 vccd1 _6164_/A sky130_fd_sc_hd__a21o_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3458_/B _4958_/A _4363_/B _3458_/A vssd1 vssd1 vccd1 vccd1 _3354_/Y sky130_fd_sc_hd__a22oi_2
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _4744_/A vssd1 vssd1 vccd1 vccd1 _5240_/B sky130_fd_sc_hd__clkbuf_4
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6205_/C _6072_/C _6072_/A _6072_/B vssd1 vssd1 vccd1 vccd1 _6073_/X sky130_fd_sc_hd__a22o_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5207_/A _5029_/B vssd1 vssd1 vccd1 vccd1 _5025_/B sky130_fd_sc_hd__nand2_4
XFILLER_38_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5926_ _5927_/C _5927_/A _5927_/B vssd1 vssd1 vccd1 vccd1 _5926_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5857_ _5850_/X _5852_/X _5848_/Y _5840_/Y vssd1 vssd1 vccd1 vccd1 _5868_/B sky130_fd_sc_hd__o211ai_4
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5788_ _5442_/C _5925_/B _5917_/C _5917_/A vssd1 vssd1 vccd1 vccd1 _5788_/Y sky130_fd_sc_hd__a22oi_4
X_4808_ _4806_/Y _4807_/Y _4639_/Y vssd1 vssd1 vccd1 vccd1 _4996_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4739_ _5397_/B vssd1 vssd1 vccd1 vccd1 _5792_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5711_ _5805_/A vssd1 vssd1 vccd1 vccd1 _5933_/C sky130_fd_sc_hd__clkbuf_2
X_3972_ _3973_/A _3973_/B _4152_/A _4011_/B vssd1 vssd1 vccd1 vccd1 _3976_/B sky130_fd_sc_hd__nand4_2
XFILLER_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5642_ _5640_/C _5640_/D _5641_/X vssd1 vssd1 vccd1 vccd1 _5643_/D sky130_fd_sc_hd__a21o_1
X_5573_ _5596_/B _5842_/A _5676_/A _5597_/A vssd1 vssd1 vccd1 vccd1 _5573_/Y sky130_fd_sc_hd__a22oi_4
X_4524_ _4524_/A vssd1 vssd1 vccd1 vccd1 _4524_/X sky130_fd_sc_hd__clkbuf_1
X_4455_ _4777_/C vssd1 vssd1 vccd1 vccd1 _5546_/A sky130_fd_sc_hd__clkbuf_4
X_3406_ _4238_/D vssd1 vssd1 vccd1 vccd1 _5663_/B sky130_fd_sc_hd__buf_4
X_4386_ _3334_/A _5808_/B _5986_/B _4186_/A vssd1 vssd1 vccd1 vccd1 _4386_/Y sky130_fd_sc_hd__a22oi_4
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3337_ _3337_/A _5905_/A _4042_/B vssd1 vssd1 vccd1 vccd1 _3487_/A sky130_fd_sc_hd__and3_1
X_6125_ _6125_/A _6127_/D vssd1 vssd1 vccd1 vccd1 _6126_/B sky130_fd_sc_hd__nand2_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6058_/B _6058_/C _6055_/X vssd1 vssd1 vccd1 vccd1 _6059_/A sky130_fd_sc_hd__a21o_1
XFILLER_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3268_ _3437_/A vssd1 vssd1 vccd1 vccd1 _3870_/A sky130_fd_sc_hd__clkbuf_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _5007_/A _5506_/A vssd1 vssd1 vccd1 vccd1 _5007_/Y sky130_fd_sc_hd__nand2_1
X_3199_ _3199_/A _3199_/B _3199_/C vssd1 vssd1 vccd1 vccd1 _3201_/A sky130_fd_sc_hd__and3_1
XFILLER_26_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5909_ _5914_/A _5914_/B _5914_/C _5998_/B vssd1 vssd1 vccd1 vccd1 _5911_/A sky130_fd_sc_hd__a22oi_1
XFILLER_14_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4240_ _4240_/A vssd1 vssd1 vccd1 vccd1 _4422_/A sky130_fd_sc_hd__clkbuf_2
X_4171_ _4010_/A _4054_/C _4010_/C _4157_/B vssd1 vssd1 vccd1 vccd1 _4171_/X sky130_fd_sc_hd__o31a_1
XFILLER_67_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3955_ input2/X vssd1 vssd1 vccd1 vccd1 _5284_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5625_ _5625_/A _5625_/B _5625_/C _5625_/D vssd1 vssd1 vccd1 vccd1 _5627_/B sky130_fd_sc_hd__nand4_1
X_3886_ _4068_/A vssd1 vssd1 vccd1 vccd1 _4460_/B sky130_fd_sc_hd__clkinv_2
X_5556_ _5561_/C vssd1 vssd1 vccd1 vccd1 _5556_/Y sky130_fd_sc_hd__clkinv_2
X_5487_ _5203_/A _5203_/B _5485_/B _5484_/A vssd1 vssd1 vccd1 vccd1 _5487_/Y sky130_fd_sc_hd__a22oi_1
X_4507_ _4681_/A _4681_/B _4516_/A _4516_/B vssd1 vssd1 vccd1 vccd1 _4514_/B sky130_fd_sc_hd__o211ai_1
XFILLER_2_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4438_ _4861_/A _4569_/A vssd1 vssd1 vccd1 vccd1 _4568_/A sky130_fd_sc_hd__nand2_4
X_4369_ _4369_/A _5539_/A vssd1 vssd1 vccd1 vccd1 _4529_/A sky130_fd_sc_hd__nand2_2
X_6108_ _6108_/A _6108_/B _6108_/C vssd1 vssd1 vccd1 vccd1 _6110_/D sky130_fd_sc_hd__nand3_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6039_ _6090_/C _5999_/B _6037_/Y _6038_/Y vssd1 vssd1 vccd1 vccd1 _6041_/B sky130_fd_sc_hd__o211ai_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_19 _5363_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3740_ _3593_/B _3488_/X _3586_/B _3586_/C vssd1 vssd1 vccd1 vccd1 _3740_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3671_ _4229_/B vssd1 vssd1 vccd1 vccd1 _5299_/B sky130_fd_sc_hd__buf_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5410_ _5701_/B vssd1 vssd1 vccd1 vccd1 _5688_/A sky130_fd_sc_hd__clkbuf_2
X_5341_ _5333_/X _5163_/X _5337_/X vssd1 vssd1 vccd1 vccd1 _5341_/Y sky130_fd_sc_hd__o21ai_1
X_5272_ _5220_/Y _5219_/X _5281_/B _5281_/A vssd1 vssd1 vccd1 vccd1 _5272_/X sky130_fd_sc_hd__o211a_1
X_4223_ _3731_/C _6233_/A _4048_/C _4177_/X vssd1 vssd1 vccd1 vccd1 _4224_/C sky130_fd_sc_hd__a31o_1
X_4154_ _4154_/A _4157_/C vssd1 vssd1 vccd1 vccd1 _4154_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4085_ _3414_/B _4935_/A _5285_/A _3551_/A vssd1 vssd1 vccd1 vccd1 _4085_/X sky130_fd_sc_hd__a22o_1
XFILLER_70_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4987_ _4988_/C _4988_/D _4971_/C vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__a21o_1
X_3938_ _3938_/A _3938_/B vssd1 vssd1 vccd1 vccd1 _3946_/A sky130_fd_sc_hd__nor2_1
X_3869_ _3280_/X _3797_/X _3787_/B _4103_/A _3868_/Y vssd1 vssd1 vccd1 vccd1 _3875_/B
+ sky130_fd_sc_hd__o221ai_2
X_5608_ _5608_/A _5608_/B _5608_/C vssd1 vssd1 vccd1 vccd1 _5608_/X sky130_fd_sc_hd__and3_1
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5539_ _5539_/A _5539_/B vssd1 vssd1 vccd1 vccd1 _5697_/A sky130_fd_sc_hd__nand2_2
XFILLER_74_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput28 b[3] vssd1 vssd1 vccd1 vccd1 _3210_/A sky130_fd_sc_hd__buf_2
Xinput17 b[10] vssd1 vssd1 vccd1 vccd1 _4252_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5890_ _5892_/B _5892_/C _5892_/A vssd1 vssd1 vccd1 vccd1 _5891_/C sky130_fd_sc_hd__a21o_1
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4910_ _4592_/B _4751_/B _4754_/A _4762_/A vssd1 vssd1 vccd1 vccd1 _4917_/A sky130_fd_sc_hd__a22o_2
X_4841_ _4842_/B _4842_/D vssd1 vssd1 vccd1 vccd1 _4841_/X sky130_fd_sc_hd__and2_1
X_4772_ _4772_/A _4924_/A _4924_/B vssd1 vssd1 vccd1 vccd1 _4801_/B sky130_fd_sc_hd__nand3_2
X_3723_ _3723_/A _3723_/B _3723_/C vssd1 vssd1 vccd1 vccd1 _3836_/A sky130_fd_sc_hd__nand3_2
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3654_ _3774_/B vssd1 vssd1 vccd1 vccd1 _4423_/A sky130_fd_sc_hd__buf_2
X_3585_ _3592_/A _3482_/A _3593_/C vssd1 vssd1 vccd1 vccd1 _3586_/A sky130_fd_sc_hd__a21bo_1
X_5324_ _5151_/Y _5153_/X _5157_/B vssd1 vssd1 vccd1 vccd1 _5325_/B sky130_fd_sc_hd__o21ai_1
X_5255_ _5244_/Y _5249_/Y _5252_/X _5268_/A _5268_/B vssd1 vssd1 vccd1 vccd1 _5256_/C
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4206_ _4384_/A vssd1 vssd1 vccd1 vccd1 _5809_/B sky130_fd_sc_hd__buf_2
X_5186_ _5173_/A _5182_/B _5185_/X vssd1 vssd1 vccd1 vccd1 _5189_/A sky130_fd_sc_hd__a21o_1
X_4137_ _4137_/A _4137_/B _4137_/C vssd1 vssd1 vccd1 vccd1 _4317_/A sky130_fd_sc_hd__nand3_2
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4068_ _4068_/A vssd1 vssd1 vccd1 vccd1 _5285_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3370_ _3368_/Y _3369_/Y _3366_/Y vssd1 vssd1 vccd1 vccd1 _3370_/X sky130_fd_sc_hd__a21o_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5040_/A _5040_/B vssd1 vssd1 vccd1 vccd1 _5041_/C sky130_fd_sc_hd__nand2_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5942_ _5942_/A _5942_/B _5942_/C vssd1 vssd1 vccd1 vccd1 _5943_/C sky130_fd_sc_hd__nand3_1
XFILLER_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5873_ _5672_/X _5685_/X _5786_/A vssd1 vssd1 vccd1 vccd1 _5873_/X sky130_fd_sc_hd__o21a_1
X_4824_ _4824_/A _4824_/B _4824_/C vssd1 vssd1 vccd1 vccd1 _4824_/Y sky130_fd_sc_hd__nand3_4
X_4755_ _4901_/B vssd1 vssd1 vccd1 vccd1 _5448_/B sky130_fd_sc_hd__buf_2
XFILLER_21_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3706_ _4855_/A _4861_/A _3758_/B _4234_/A vssd1 vssd1 vccd1 vccd1 _3754_/B sky130_fd_sc_hd__nand4_1
X_4686_ _4686_/A _4686_/B vssd1 vssd1 vccd1 vccd1 _4686_/Y sky130_fd_sc_hd__xnor2_4
X_3637_ _3625_/Y _3691_/A _3635_/X _3636_/Y vssd1 vssd1 vccd1 vccd1 _3720_/A sky130_fd_sc_hd__o2bb2ai_2
X_3568_ _3568_/A vssd1 vssd1 vccd1 vccd1 _3703_/B sky130_fd_sc_hd__clkbuf_2
X_5307_ _5307_/A _5307_/B _5307_/C vssd1 vssd1 vccd1 vccd1 _5321_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6287_ _6287_/A _6292_/B vssd1 vssd1 vccd1 vccd1 _6289_/A sky130_fd_sc_hd__nand2_1
X_3499_ _3514_/A _5578_/A _3508_/D _3504_/A vssd1 vssd1 vccd1 vccd1 _3509_/A sky130_fd_sc_hd__a22o_1
X_5238_ _5238_/A vssd1 vssd1 vccd1 vccd1 _5677_/A sky130_fd_sc_hd__buf_2
X_5169_ _5175_/A _5175_/B vssd1 vssd1 vccd1 vccd1 _5170_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4540_ _4540_/A _4540_/B _4708_/C _5299_/D vssd1 vssd1 vccd1 vccd1 _4540_/Y sky130_fd_sc_hd__nand4_1
X_4471_ _4464_/X _4266_/Y _4270_/Y _4298_/D _4294_/C vssd1 vssd1 vccd1 vccd1 _4478_/A
+ sky130_fd_sc_hd__a32o_1
X_6210_ _6178_/B _6183_/A _6227_/A vssd1 vssd1 vccd1 vccd1 _6212_/A sky130_fd_sc_hd__o21a_1
X_3422_ _4884_/A vssd1 vssd1 vccd1 vccd1 _4236_/A sky130_fd_sc_hd__clkbuf_4
X_6141_ _6138_/A _6138_/B _6131_/X _6140_/Y vssd1 vssd1 vccd1 vccd1 _6143_/B sky130_fd_sc_hd__o22ai_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _4369_/A vssd1 vssd1 vccd1 vccd1 _4363_/B sky130_fd_sc_hd__buf_2
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3908_/A vssd1 vssd1 vccd1 vccd1 _4744_/A sky130_fd_sc_hd__buf_2
X_6072_ _6072_/A _6072_/B _6072_/C vssd1 vssd1 vccd1 vccd1 _6072_/Y sky130_fd_sc_hd__nand3_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5021_/A _4986_/X _5021_/C vssd1 vssd1 vccd1 vccd1 _5172_/A sky130_fd_sc_hd__o21ai_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5925_ _5925_/A _5925_/B vssd1 vssd1 vccd1 vccd1 _5927_/B sky130_fd_sc_hd__and2_1
X_5856_ _5840_/Y _5848_/Y _5855_/X vssd1 vssd1 vccd1 vccd1 _5868_/A sky130_fd_sc_hd__a21o_2
X_4807_ _4639_/A _4639_/B _4639_/C vssd1 vssd1 vccd1 vccd1 _4807_/Y sky130_fd_sc_hd__a21oi_1
X_5787_ _5860_/A _5786_/Y _5747_/Y _5756_/Y vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__o22ai_2
XFILLER_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4738_ _4738_/A _5059_/A vssd1 vssd1 vccd1 vccd1 _4853_/A sky130_fd_sc_hd__nand2_1
X_4669_ _4669_/A vssd1 vssd1 vccd1 vccd1 _4669_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3971_ _4010_/A _4052_/A _4010_/C vssd1 vssd1 vccd1 vccd1 _4011_/B sky130_fd_sc_hd__o21ai_1
X_5710_ _5726_/A vssd1 vssd1 vccd1 vccd1 _5728_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5641_ _4417_/X _4674_/X _5438_/Y _5640_/A vssd1 vssd1 vccd1 vccd1 _5641_/X sky130_fd_sc_hd__o31a_1
X_5572_ _5658_/A vssd1 vssd1 vccd1 vccd1 _5842_/A sky130_fd_sc_hd__buf_2
X_4523_ _4513_/X _4518_/X _4523_/S vssd1 vssd1 vccd1 vccd1 _4524_/A sky130_fd_sc_hd__mux2_4
X_4454_ _5374_/A _4454_/B _5223_/A _4761_/B vssd1 vssd1 vccd1 vccd1 _4456_/B sky130_fd_sc_hd__nand4_1
X_4385_ _5434_/D vssd1 vssd1 vccd1 vccd1 _5986_/B sky130_fd_sc_hd__clkbuf_4
X_3405_ _4906_/A vssd1 vssd1 vccd1 vccd1 _4238_/D sky130_fd_sc_hd__clkbuf_4
X_6124_ _6124_/A _6124_/B vssd1 vssd1 vccd1 vccd1 _6236_/C sky130_fd_sc_hd__nand2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ _3731_/C _5905_/A _3337_/A vssd1 vssd1 vccd1 vccd1 _3389_/A sky130_fd_sc_hd__a21oi_1
X_6055_ _6058_/A _5969_/C _5969_/B vssd1 vssd1 vccd1 vccd1 _6055_/X sky130_fd_sc_hd__a21bo_1
XFILLER_85_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5006_ _5006_/A _5348_/D vssd1 vssd1 vccd1 vccd1 _5006_/Y sky130_fd_sc_hd__nand2_1
X_3267_ _3500_/A vssd1 vssd1 vccd1 vccd1 _4547_/A sky130_fd_sc_hd__buf_4
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3198_ _3966_/A _3310_/C vssd1 vssd1 vccd1 vccd1 _3199_/C sky130_fd_sc_hd__nand2_1
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5908_ _5914_/D vssd1 vssd1 vccd1 vccd1 _5998_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5839_ _5662_/B _6096_/A _5852_/C _6170_/C _5914_/A vssd1 vssd1 vccd1 vccd1 _5840_/C
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_5_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4170_ _4008_/X _4012_/Y _4138_/Y _4145_/Y vssd1 vssd1 vccd1 vccd1 _4170_/X sky130_fd_sc_hd__o211a_1
XFILLER_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3954_ _5541_/A vssd1 vssd1 vccd1 vccd1 _5919_/A sky130_fd_sc_hd__clkbuf_4
X_3885_ _3650_/Y _3891_/A _3758_/Y _3760_/Y vssd1 vssd1 vccd1 vccd1 _4096_/A sky130_fd_sc_hd__o22a_1
XFILLER_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5624_ _5624_/A _5624_/B vssd1 vssd1 vccd1 vccd1 _5627_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5555_ _5555_/A _5555_/B _5555_/C vssd1 vssd1 vccd1 vccd1 _5561_/C sky130_fd_sc_hd__nand3_4
X_5486_ _5327_/Y _5495_/A _5329_/X vssd1 vssd1 vccd1 vccd1 _5486_/Y sky130_fd_sc_hd__o21ai_1
X_4506_ _4506_/A _4506_/B _4506_/C vssd1 vssd1 vccd1 vccd1 _4516_/B sky130_fd_sc_hd__nand3_1
X_4437_ _4435_/Y _4436_/Y _4277_/B vssd1 vssd1 vccd1 vccd1 _4601_/B sky130_fd_sc_hd__o21ai_2
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6107_ _6108_/A _6108_/B _6108_/C vssd1 vssd1 vccd1 vccd1 _6159_/A sky130_fd_sc_hd__a21o_1
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ _4958_/B _5696_/A _5701_/A _4547_/A vssd1 vssd1 vccd1 vccd1 _4368_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4299_ _4298_/A _4298_/B _4298_/C _4298_/D vssd1 vssd1 vccd1 vccd1 _4299_/X sky130_fd_sc_hd__a22o_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _5207_/A vssd1 vssd1 vccd1 vccd1 _5209_/A sky130_fd_sc_hd__clkbuf_4
X_6038_ _6024_/Y _6022_/Y _6034_/B _6030_/Y vssd1 vssd1 vccd1 vccd1 _6038_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3670_ _5603_/A _3669_/X _3656_/A vssd1 vssd1 vccd1 vccd1 _3708_/B sky130_fd_sc_hd__o21ai_1
X_5340_ _5323_/B _5323_/C _5323_/A vssd1 vssd1 vccd1 vccd1 _5340_/Y sky130_fd_sc_hd__a21oi_2
X_5271_ _5271_/A vssd1 vssd1 vccd1 vccd1 _5281_/B sky130_fd_sc_hd__buf_2
X_4222_ _6170_/A vssd1 vssd1 vccd1 vccd1 _6233_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4153_ _4157_/A _4157_/B vssd1 vssd1 vccd1 vccd1 _4154_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4084_ _4877_/B _4234_/A vssd1 vssd1 vccd1 vccd1 _4254_/A sky130_fd_sc_hd__nand2_2
XFILLER_55_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4986_ _4927_/Y _4973_/Y _4979_/Y _4985_/Y vssd1 vssd1 vccd1 vccd1 _4986_/X sky130_fd_sc_hd__o211a_1
X_3937_ _3945_/A _3984_/C vssd1 vssd1 vccd1 vccd1 _3939_/A sky130_fd_sc_hd__nand2_1
X_3868_ _3868_/A _3868_/B vssd1 vssd1 vccd1 vccd1 _3868_/Y sky130_fd_sc_hd__nand2_2
X_5607_ _5590_/Y _5686_/A _5686_/B _5609_/B vssd1 vssd1 vccd1 vccd1 _5611_/A sky130_fd_sc_hd__nand4b_4
X_3799_ _3799_/A _3799_/B _3799_/C vssd1 vssd1 vccd1 vccd1 _3799_/Y sky130_fd_sc_hd__nand3_2
X_5538_ _5538_/A vssd1 vssd1 vccd1 vccd1 _5538_/X sky130_fd_sc_hd__buf_2
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5469_ _4907_/X _5025_/B _3634_/X _4287_/B vssd1 vssd1 vccd1 vccd1 _5469_/X sky130_fd_sc_hd__a211o_1
XFILLER_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 b[11] vssd1 vssd1 vccd1 vccd1 _4260_/A sky130_fd_sc_hd__clkbuf_1
Xinput29 b[4] vssd1 vssd1 vccd1 vccd1 _3356_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4840_ _4508_/Y _4525_/X _4672_/Y _4676_/X vssd1 vssd1 vccd1 vccd1 _4840_/X sky130_fd_sc_hd__o211a_1
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _4742_/X _4749_/Y _4762_/X _4763_/Y vssd1 vssd1 vccd1 vccd1 _4924_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_9_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3722_ _3561_/A _3702_/A _3702_/B _3568_/A _3703_/A vssd1 vssd1 vccd1 vccd1 _3723_/C
+ sky130_fd_sc_hd__a32oi_2
X_3653_ _3646_/Y _3650_/Y _3747_/A _3530_/B vssd1 vssd1 vccd1 vccd1 _3656_/A sky130_fd_sc_hd__o2bb2ai_1
X_5323_ _5323_/A _5323_/B _5323_/C vssd1 vssd1 vccd1 vccd1 _5337_/A sky130_fd_sc_hd__nand3_1
X_3584_ _3584_/A _3584_/B _3584_/C vssd1 vssd1 vccd1 vccd1 _3593_/C sky130_fd_sc_hd__nand3_2
XFILLER_87_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5254_ _5420_/A _5254_/B vssd1 vssd1 vccd1 vccd1 _5256_/B sky130_fd_sc_hd__nand2_1
X_5185_ _4943_/C _5352_/A _5006_/A _4958_/X vssd1 vssd1 vccd1 vccd1 _5185_/X sky130_fd_sc_hd__a31o_1
X_4205_ _5808_/B vssd1 vssd1 vccd1 vccd1 _6077_/A sky130_fd_sc_hd__buf_4
X_4136_ _4134_/Y _4135_/X _4124_/C _4124_/A vssd1 vssd1 vccd1 vccd1 _4137_/C sky130_fd_sc_hd__o211ai_4
XFILLER_56_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4067_ _4067_/A _5240_/A _5284_/C _5212_/B vssd1 vssd1 vccd1 vccd1 _4067_/Y sky130_fd_sc_hd__nand4_4
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4969_ _4722_/A _4722_/B _4721_/X vssd1 vssd1 vccd1 vccd1 _4971_/C sky130_fd_sc_hd__a21oi_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5941_ _5942_/C _5937_/A _5935_/A _5935_/B vssd1 vssd1 vccd1 vccd1 _5943_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5872_ _5872_/A _5872_/B _5872_/C vssd1 vssd1 vccd1 vccd1 _5872_/Y sky130_fd_sc_hd__nand3_2
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4823_ _4661_/A _4661_/B _4661_/C _4663_/A _4669_/Y vssd1 vssd1 vccd1 vccd1 _4824_/C
+ sky130_fd_sc_hd__a32oi_4
X_4754_ _4754_/A vssd1 vssd1 vccd1 vccd1 _4890_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3705_ _3705_/A _3705_/B _3705_/C vssd1 vssd1 vccd1 vccd1 _3835_/A sky130_fd_sc_hd__nand3_2
X_4685_ _4523_/S _4513_/X _4842_/B vssd1 vssd1 vccd1 vccd1 _4686_/B sky130_fd_sc_hd__o21ai_2
X_3636_ _4827_/A _5905_/A _5994_/A _3829_/B vssd1 vssd1 vccd1 vccd1 _3636_/Y sky130_fd_sc_hd__a22oi_2
X_3567_ _3567_/A _3567_/B _3567_/C vssd1 vssd1 vccd1 vccd1 _3568_/A sky130_fd_sc_hd__nand3_1
X_6286_ _6286_/A _6285_/A vssd1 vssd1 vccd1 vccd1 _6292_/B sky130_fd_sc_hd__or2b_1
X_5306_ _5032_/B _5032_/C _5032_/A _5309_/A _5309_/B vssd1 vssd1 vccd1 vccd1 _5307_/C
+ sky130_fd_sc_hd__a32oi_1
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3498_ _3498_/A _3498_/B vssd1 vssd1 vccd1 vccd1 _3504_/A sky130_fd_sc_hd__nand2_1
X_5237_ _5237_/A vssd1 vssd1 vccd1 vccd1 _5831_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5168_ _4968_/A _4968_/B _4968_/C _4971_/C vssd1 vssd1 vccd1 vccd1 _5175_/B sky130_fd_sc_hd__a31o_1
X_5099_ _4917_/B _4917_/C _4917_/A vssd1 vssd1 vccd1 vccd1 _5099_/Y sky130_fd_sc_hd__a21oi_2
X_4119_ _4135_/C vssd1 vssd1 vccd1 vccd1 _4220_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4470_ _4308_/B _4303_/Y _4296_/A vssd1 vssd1 vccd1 vccd1 _4470_/Y sky130_fd_sc_hd__a21boi_1
X_3421_ _4540_/B _5251_/A _4708_/B _5373_/A vssd1 vssd1 vccd1 vccd1 _3421_/Y sky130_fd_sc_hd__nand4_2
X_6140_ _6132_/Y _6129_/Y _6130_/X vssd1 vssd1 vccd1 vccd1 _6140_/Y sky130_fd_sc_hd__a21oi_1
X_3352_ _3500_/A vssd1 vssd1 vccd1 vccd1 _4958_/A sky130_fd_sc_hd__clkbuf_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6071_ _6071_/A vssd1 vssd1 vccd1 vccd1 _6072_/C sky130_fd_sc_hd__buf_2
X_3283_ _3533_/B _4369_/A vssd1 vssd1 vccd1 vccd1 _3342_/A sky130_fd_sc_hd__nand2_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5019_/Y _5005_/Y _5020_/Y _5021_/X vssd1 vssd1 vccd1 vccd1 _5184_/A sky130_fd_sc_hd__o2bb2a_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5924_ _6025_/A _6025_/B _6025_/C vssd1 vssd1 vccd1 vccd1 _5942_/C sky130_fd_sc_hd__nand3_2
XFILLER_53_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5855_ _6096_/C _5852_/A _5825_/D _5850_/X vssd1 vssd1 vccd1 vccd1 _5855_/X sky130_fd_sc_hd__a31o_1
XFILLER_61_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4806_ _4806_/A _4817_/B vssd1 vssd1 vccd1 vccd1 _4806_/Y sky130_fd_sc_hd__nand2_1
X_5786_ _5786_/A _5786_/B vssd1 vssd1 vccd1 vccd1 _5786_/Y sky130_fd_sc_hd__nand2_1
X_4737_ _4573_/A _4579_/Y _4576_/C vssd1 vssd1 vccd1 vccd1 _4741_/B sky130_fd_sc_hd__o21ai_1
X_4668_ _4400_/C _4395_/Y _4400_/A _4663_/B _4663_/A vssd1 vssd1 vccd1 vccd1 _4671_/B
+ sky130_fd_sc_hd__o2111ai_4
X_3619_ _5029_/A vssd1 vssd1 vccd1 vccd1 _5399_/A sky130_fd_sc_hd__buf_4
X_4599_ _4599_/A _4599_/B vssd1 vssd1 vccd1 vccd1 _4607_/A sky130_fd_sc_hd__nand2_1
X_6269_ _6224_/B _6223_/X _6274_/A _6197_/B vssd1 vssd1 vccd1 vccd1 _6271_/A sky130_fd_sc_hd__o22ai_1
XFILLER_0_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3970_ _4010_/A _4052_/A _4010_/C vssd1 vssd1 vccd1 vccd1 _4152_/A sky130_fd_sc_hd__or3_2
XFILLER_43_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5640_ _5640_/A _5640_/B _5640_/C _5640_/D vssd1 vssd1 vccd1 vccd1 _5643_/C sky130_fd_sc_hd__nand4_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5571_ _5594_/A _6002_/B vssd1 vssd1 vccd1 vccd1 _5571_/Y sky130_fd_sc_hd__nand2_1
X_4522_ _4519_/X _4520_/Y _4521_/Y _4164_/Y vssd1 vssd1 vccd1 vccd1 _4523_/S sky130_fd_sc_hd__a22oi_4
XFILLER_7_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4453_ _4454_/B _5223_/A _4761_/B _5374_/A vssd1 vssd1 vccd1 vccd1 _4453_/Y sky130_fd_sc_hd__a22oi_4
X_3404_ _3473_/A _5211_/A vssd1 vssd1 vccd1 vccd1 _3498_/A sky130_fd_sc_hd__nand2_2
X_4384_ _4384_/A vssd1 vssd1 vccd1 vccd1 _5434_/D sky130_fd_sc_hd__clkbuf_2
X_6123_ _6101_/A _6101_/B _6104_/A vssd1 vssd1 vccd1 vccd1 _6123_/X sky130_fd_sc_hd__a21o_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3335_ _3265_/A _5678_/B _3521_/A _3334_/X vssd1 vssd1 vccd1 vccd1 _3337_/A sky130_fd_sc_hd__a31o_1
X_6054_ _6054_/A _6054_/B vssd1 vssd1 vccd1 vccd1 _6058_/C sky130_fd_sc_hd__nand2_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _3356_/A vssd1 vssd1 vccd1 vccd1 _3500_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5005_ _5005_/A _5005_/B _5005_/C vssd1 vssd1 vccd1 vccd1 _5005_/Y sky130_fd_sc_hd__nand3_4
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3197_ _5597_/A vssd1 vssd1 vccd1 vccd1 _3310_/C sky130_fd_sc_hd__buf_2
XFILLER_66_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5907_ _5907_/A _5998_/A _6096_/C _6203_/C vssd1 vssd1 vccd1 vccd1 _5914_/D sky130_fd_sc_hd__nand4_2
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5838_ _5846_/A vssd1 vssd1 vccd1 vccd1 _5914_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5769_ _5535_/X _5352_/A _4621_/C _5532_/X vssd1 vssd1 vccd1 vccd1 _5781_/B sky130_fd_sc_hd__a31o_1
XFILLER_14_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3953_ _5123_/B vssd1 vssd1 vccd1 vccd1 _5541_/A sky130_fd_sc_hd__clkbuf_4
X_3884_ _4430_/A _4065_/A vssd1 vssd1 vccd1 vccd1 _3891_/A sky130_fd_sc_hd__nand2_2
X_5623_ _5623_/A _5623_/B vssd1 vssd1 vccd1 vccd1 _5624_/B sky130_fd_sc_hd__nand2_1
X_5554_ _5554_/A _5554_/B vssd1 vssd1 vccd1 vccd1 _5555_/C sky130_fd_sc_hd__nand2_1
X_5485_ _5485_/A _5485_/B vssd1 vssd1 vccd1 vccd1 _5485_/Y sky130_fd_sc_hd__nand2_1
X_4505_ _4506_/C _4506_/B _4506_/A vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__a21o_1
X_4436_ _3533_/B _4884_/B _4753_/D _3533_/A vssd1 vssd1 vccd1 vccd1 _4436_/Y sky130_fd_sc_hd__a22oi_4
X_4367_ _4363_/Y _4365_/Y _4366_/Y vssd1 vssd1 vccd1 vccd1 _4367_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6106_ _6047_/A _6105_/Y _6047_/B vssd1 vssd1 vccd1 vccd1 _6108_/C sky130_fd_sc_hd__a21bo_1
XFILLER_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3318_ _4901_/A vssd1 vssd1 vccd1 vccd1 _5207_/A sky130_fd_sc_hd__buf_2
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4298_ _4298_/A _4298_/B _4298_/C _4298_/D vssd1 vssd1 vccd1 vccd1 _4298_/Y sky130_fd_sc_hd__nand4_2
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6037_ _6037_/A _6037_/B vssd1 vssd1 vccd1 vccd1 _6037_/Y sky130_fd_sc_hd__nand2_1
X_3249_ _3256_/A vssd1 vssd1 vccd1 vccd1 _4193_/A sky130_fd_sc_hd__buf_2
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5270_ _5221_/X _5226_/X _5490_/A _5431_/A vssd1 vssd1 vccd1 vccd1 _5277_/B sky130_fd_sc_hd__o211ai_2
X_4221_ _5808_/B vssd1 vssd1 vccd1 vccd1 _6170_/A sky130_fd_sc_hd__clkbuf_2
X_4152_ _4152_/A _4157_/A _4157_/B vssd1 vssd1 vccd1 vccd1 _4152_/Y sky130_fd_sc_hd__nand3_1
XFILLER_95_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4083_ _4284_/A _4284_/B _4284_/C vssd1 vssd1 vccd1 vccd1 _4100_/B sky130_fd_sc_hd__nand3_4
XFILLER_95_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4985_ _4985_/A _4985_/B vssd1 vssd1 vccd1 vccd1 _4985_/Y sky130_fd_sc_hd__nand2_2
X_3936_ _3936_/A vssd1 vssd1 vccd1 vccd1 _3984_/C sky130_fd_sc_hd__clkbuf_1
X_3867_ _3867_/A _5655_/A vssd1 vssd1 vccd1 vccd1 _3868_/B sky130_fd_sc_hd__nand2_1
X_3798_ _3468_/A _3797_/X _3791_/A _3791_/B vssd1 vssd1 vccd1 vccd1 _3799_/C sky130_fd_sc_hd__o211ai_1
X_5606_ _5603_/X _5612_/A _5604_/X _5605_/Y vssd1 vssd1 vccd1 vccd1 _5609_/B sky130_fd_sc_hd__o2bb2ai_4
X_5537_ _5694_/A _5694_/B vssd1 vssd1 vccd1 vccd1 _5550_/A sky130_fd_sc_hd__nand2_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5468_ _5640_/B _5468_/B _5468_/C _5468_/D vssd1 vssd1 vccd1 vccd1 _5471_/B sky130_fd_sc_hd__nand4_1
X_4419_ _4405_/Y _4415_/X _4416_/Y _4418_/Y vssd1 vssd1 vccd1 vccd1 _4420_/A sky130_fd_sc_hd__o211ai_1
X_5399_ _5399_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _5399_/Y sky130_fd_sc_hd__nand2_4
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput19 b[12] vssd1 vssd1 vccd1 vccd1 _4078_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4770_ _4757_/Y _4758_/X _4768_/Y _4769_/Y _4742_/X vssd1 vssd1 vccd1 vccd1 _4924_/A
+ sky130_fd_sc_hd__o221ai_4
X_3721_ _3720_/A _3720_/B _3720_/C _3720_/D vssd1 vssd1 vccd1 vccd1 _3723_/B sky130_fd_sc_hd__a22o_1
X_3652_ _4430_/A _4068_/A vssd1 vssd1 vccd1 vccd1 _3747_/A sky130_fd_sc_hd__nand2_2
X_3583_ _3593_/B _3488_/X _3586_/B _3586_/C vssd1 vssd1 vccd1 vccd1 _3857_/A sky130_fd_sc_hd__a22o_1
X_5322_ _5320_/Y _5321_/X _5277_/Y _5283_/Y vssd1 vssd1 vccd1 vccd1 _5323_/C sky130_fd_sc_hd__o211ai_2
X_5253_ _5244_/Y _5249_/Y _5252_/X vssd1 vssd1 vccd1 vccd1 _5254_/B sky130_fd_sc_hd__o21ai_1
X_5184_ _5184_/A _5184_/B _5184_/C vssd1 vssd1 vccd1 vccd1 _5517_/A sky130_fd_sc_hd__nand3_2
X_4204_ _4708_/C vssd1 vssd1 vccd1 vccd1 _5808_/B sky130_fd_sc_hd__buf_2
XFILLER_68_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4135_ _4127_/C _4135_/B _4135_/C vssd1 vssd1 vccd1 vccd1 _4135_/X sky130_fd_sc_hd__and3b_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4066_ _4906_/B vssd1 vssd1 vccd1 vccd1 _5212_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_71_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4968_ _4968_/A _4968_/B _4968_/C vssd1 vssd1 vccd1 vccd1 _4988_/D sky130_fd_sc_hd__nand3_1
X_4899_ _4981_/B _4981_/C vssd1 vssd1 vccd1 vccd1 _4921_/A sky130_fd_sc_hd__nand2_1
X_3919_ _3927_/A _3912_/A _3917_/X _3918_/X vssd1 vssd1 vccd1 vccd1 _3920_/C sky130_fd_sc_hd__o2bb2ai_1
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5940_ _5940_/A _5940_/B _5940_/C vssd1 vssd1 vccd1 vccd1 _5940_/Y sky130_fd_sc_hd__nand3_2
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5871_ _5865_/X _5866_/Y _5870_/Y vssd1 vssd1 vccd1 vccd1 _5872_/C sky130_fd_sc_hd__o21ai_1
XFILLER_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4822_ _4822_/A _4822_/B _4822_/C vssd1 vssd1 vccd1 vccd1 _4824_/B sky130_fd_sc_hd__nand3_1
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4753_ _5066_/A _5068_/B _4884_/B _4753_/D vssd1 vssd1 vccd1 vccd1 _4754_/A sky130_fd_sc_hd__nand4_2
X_3704_ _3567_/B _3702_/Y _3703_/Y vssd1 vssd1 vccd1 vccd1 _3705_/C sky130_fd_sc_hd__o21ai_1
X_4684_ _4842_/C _4842_/D vssd1 vssd1 vccd1 vccd1 _4686_/A sky130_fd_sc_hd__nand2_2
X_3635_ _3186_/X _3634_/X _3498_/A _3498_/B vssd1 vssd1 vccd1 vccd1 _3635_/X sky130_fd_sc_hd__o22a_1
X_3566_ _3564_/X _3565_/Y _3560_/B _3558_/A vssd1 vssd1 vccd1 vccd1 _3567_/C sky130_fd_sc_hd__o211ai_1
X_6285_ _6285_/A _6286_/A vssd1 vssd1 vccd1 vccd1 _6287_/A sky130_fd_sc_hd__or2b_1
X_5305_ _5289_/Y _5293_/Y _5303_/A _5303_/B _5297_/Y vssd1 vssd1 vccd1 vccd1 _5307_/B
+ sky130_fd_sc_hd__o221ai_1
X_3497_ _4714_/A _5655_/A vssd1 vssd1 vccd1 vccd1 _3498_/B sky130_fd_sc_hd__nand2_1
XFILLER_88_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5236_ _5236_/A _5236_/B vssd1 vssd1 vccd1 vccd1 _5268_/A sky130_fd_sc_hd__nand2_2
X_5167_ _5171_/C _5171_/D vssd1 vssd1 vccd1 vccd1 _5176_/A sky130_fd_sc_hd__nand2_1
X_5098_ _5278_/A vssd1 vssd1 vccd1 vccd1 _5098_/Y sky130_fd_sc_hd__inv_2
X_4118_ _4135_/C _4211_/A _4127_/C vssd1 vssd1 vccd1 vccd1 _4122_/A sky130_fd_sc_hd__a21o_1
XFILLER_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4049_ _4048_/B _4048_/C _4047_/A vssd1 vssd1 vccd1 vccd1 _4049_/X sky130_fd_sc_hd__a21o_1
XFILLER_71_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3420_ _3468_/A _3474_/A _3368_/B _3552_/A _3419_/Y vssd1 vssd1 vccd1 vccd1 _3465_/A
+ sky130_fd_sc_hd__o221ai_4
X_3351_ _3358_/D _3440_/A _4747_/A _3350_/Y vssd1 vssd1 vccd1 vccd1 _3359_/A sky130_fd_sc_hd__o2bb2ai_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3437_/A vssd1 vssd1 vccd1 vccd1 _4369_/A sky130_fd_sc_hd__buf_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6067_/Y _6068_/X _6069_/Y vssd1 vssd1 vccd1 vccd1 _6089_/C sky130_fd_sc_hd__o21bai_4
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5021_/A _5021_/B _5021_/C vssd1 vssd1 vccd1 vccd1 _5021_/X sky130_fd_sc_hd__and3_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5923_ _5789_/Y _5788_/Y _5794_/Y vssd1 vssd1 vccd1 vccd1 _6025_/C sky130_fd_sc_hd__o21ai_1
X_5854_ _5867_/A _6236_/B _5849_/Y _5853_/X vssd1 vssd1 vccd1 vccd1 _5860_/B sky130_fd_sc_hd__o22ai_4
XFILLER_21_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4805_ _4809_/A _4809_/B _4814_/A vssd1 vssd1 vccd1 vccd1 _4996_/A sky130_fd_sc_hd__o21ai_1
X_5785_ _5673_/Y _5675_/X _5741_/Y vssd1 vssd1 vccd1 vccd1 _5860_/A sky130_fd_sc_hd__o21a_1
XFILLER_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4736_ _4746_/A _4746_/B _3441_/X _6171_/A vssd1 vssd1 vccd1 vccd1 _4741_/A sky130_fd_sc_hd__o2bb2ai_1
X_4667_ _4502_/C _4502_/A _4526_/Y vssd1 vssd1 vccd1 vccd1 _4671_/A sky130_fd_sc_hd__a21oi_4
X_3618_ _4906_/A vssd1 vssd1 vccd1 vccd1 _5029_/A sky130_fd_sc_hd__buf_2
X_4598_ _4598_/A vssd1 vssd1 vccd1 vccd1 _4599_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3549_ _3565_/A _3549_/B _3565_/B vssd1 vssd1 vccd1 vccd1 _3558_/B sky130_fd_sc_hd__nand3_2
XFILLER_95_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6268_ _6248_/A _6251_/A _6267_/Y vssd1 vssd1 vccd1 vccd1 _6273_/A sky130_fd_sc_hd__o21bai_1
XFILLER_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5219_ _3512_/X _4287_/B _4903_/B _5208_/A vssd1 vssd1 vccd1 vccd1 _5219_/X sky130_fd_sc_hd__o22a_1
X_6199_ _6199_/A _6240_/C vssd1 vssd1 vccd1 vccd1 _6257_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5570_ _5570_/A vssd1 vssd1 vccd1 vccd1 _6002_/B sky130_fd_sc_hd__clkbuf_4
X_4521_ _4340_/A _4340_/B _4338_/Y vssd1 vssd1 vccd1 vccd1 _4521_/Y sky130_fd_sc_hd__a21oi_1
X_4452_ _5286_/B vssd1 vssd1 vccd1 vccd1 _5223_/A sky130_fd_sc_hd__buf_2
X_3403_ _4906_/A vssd1 vssd1 vccd1 vccd1 _5211_/A sky130_fd_sc_hd__buf_4
X_4383_ _4237_/X _4241_/X _4381_/Y _4247_/A _4382_/X vssd1 vssd1 vccd1 vccd1 _4397_/B
+ sky130_fd_sc_hd__a32oi_4
X_6122_ _6084_/A _6084_/B _6081_/A vssd1 vssd1 vccd1 vccd1 _6156_/A sky130_fd_sc_hd__o21ai_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _3334_/A _4542_/A _5596_/A _5596_/B vssd1 vssd1 vccd1 vccd1 _3334_/X sky130_fd_sc_hd__and4_1
X_6053_ _5811_/A _6017_/A _5987_/Y vssd1 vssd1 vccd1 vccd1 _6054_/B sky130_fd_sc_hd__o21a_1
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3265_/A _5263_/C _4390_/A _3265_/D vssd1 vssd1 vccd1 vccd1 _3306_/B sky130_fd_sc_hd__nand4_2
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5021_/C _5004_/B _5021_/B vssd1 vssd1 vccd1 vccd1 _5005_/C sky130_fd_sc_hd__nand3_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3196_ _5066_/A vssd1 vssd1 vccd1 vccd1 _5597_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5906_ _6096_/C _6203_/C _5907_/A _5998_/A vssd1 vssd1 vccd1 vccd1 _5914_/C sky130_fd_sc_hd__a22o_1
X_5837_ _6001_/C vssd1 vssd1 vccd1 vccd1 _6170_/C sky130_fd_sc_hd__clkbuf_2
X_5768_ _5763_/Y _5768_/B _5768_/C vssd1 vssd1 vccd1 vccd1 _5782_/A sky130_fd_sc_hd__nand3b_1
X_4719_ _4628_/A _4628_/B _4628_/C _4635_/A _4635_/C vssd1 vssd1 vccd1 vccd1 _4719_/Y
+ sky130_fd_sc_hd__a32oi_4
X_5699_ _5809_/A _4186_/B _5799_/A _5698_/Y vssd1 vssd1 vccd1 vccd1 _5703_/A sky130_fd_sc_hd__a22o_1
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3952_ _3952_/A vssd1 vssd1 vccd1 vccd1 _5123_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3883_ _3780_/X _3764_/A _3810_/Y vssd1 vssd1 vccd1 vccd1 _3920_/A sky130_fd_sc_hd__a21oi_1
X_5622_ _5622_/A _5622_/B _5622_/C vssd1 vssd1 vccd1 vccd1 _5634_/C sky130_fd_sc_hd__nand3_2
X_5553_ _5805_/A _5553_/B vssd1 vssd1 vccd1 vccd1 _5554_/B sky130_fd_sc_hd__and2_1
X_4504_ _4503_/Y _4331_/B _4333_/B vssd1 vssd1 vccd1 vccd1 _4506_/A sky130_fd_sc_hd__o21ai_1
X_5484_ _5484_/A vssd1 vssd1 vccd1 vccd1 _5484_/Y sky130_fd_sc_hd__inv_2
X_4435_ _5231_/A _5206_/A vssd1 vssd1 vccd1 vccd1 _4435_/Y sky130_fd_sc_hd__nand2_1
X_4366_ _4366_/A _5553_/B vssd1 vssd1 vccd1 vccd1 _4366_/Y sky130_fd_sc_hd__nand2_2
XFILLER_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6105_ _6105_/A vssd1 vssd1 vccd1 vccd1 _6105_/Y sky130_fd_sc_hd__inv_2
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ _3317_/A _3317_/B vssd1 vssd1 vccd1 vccd1 _3317_/Y sky130_fd_sc_hd__nor2_4
XFILLER_86_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4297_ _4249_/Y _4250_/X _4281_/X _4291_/Y _4308_/A vssd1 vssd1 vccd1 vccd1 _4297_/Y
+ sky130_fd_sc_hd__o221ai_4
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6041_/A vssd1 vssd1 vccd1 vccd1 _6101_/A sky130_fd_sc_hd__clkbuf_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _3240_/C _3240_/A _3240_/B vssd1 vssd1 vccd1 vccd1 _3302_/A sky130_fd_sc_hd__a21bo_1
X_3179_ _3218_/A _3791_/C _3179_/C _4941_/A vssd1 vssd1 vccd1 vccd1 _3184_/D sky130_fd_sc_hd__nand4_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4220_ _4220_/A _4220_/B _4220_/C _4220_/D vssd1 vssd1 vccd1 vccd1 _4225_/A sky130_fd_sc_hd__nand4_1
X_4151_ _4151_/A vssd1 vssd1 vccd1 vccd1 _4157_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4082_ _3891_/A _4064_/X _4067_/Y _4069_/Y vssd1 vssd1 vccd1 vccd1 _4284_/C sky130_fd_sc_hd__a22oi_4
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4984_ _4984_/A _4984_/B vssd1 vssd1 vccd1 vccd1 _4985_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3935_ _3930_/Y _3931_/Y _3822_/C _3934_/Y vssd1 vssd1 vccd1 vccd1 _3985_/A sky130_fd_sc_hd__a22oi_4
XFILLER_23_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3866_ _3866_/A _4904_/B vssd1 vssd1 vccd1 vccd1 _3868_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5605_ _5604_/B _5661_/A _5604_/A vssd1 vssd1 vccd1 vccd1 _5605_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3797_ _5034_/A vssd1 vssd1 vccd1 vccd1 _3797_/X sky130_fd_sc_hd__clkbuf_4
X_5536_ _3669_/X _4711_/C _5437_/B _5534_/Y _5535_/X vssd1 vssd1 vccd1 vccd1 _5694_/B
+ sky130_fd_sc_hd__o221ai_4
X_5467_ _5640_/B _5468_/B _5468_/C _5468_/D vssd1 vssd1 vccd1 vccd1 _5471_/A sky130_fd_sc_hd__a22o_1
X_4418_ _4410_/Y _4630_/A _4417_/X _3634_/A vssd1 vssd1 vccd1 vccd1 _4418_/Y sky130_fd_sc_hd__o2bb2ai_1
X_5398_ _5403_/B vssd1 vssd1 vccd1 vccd1 _5674_/A sky130_fd_sc_hd__clkbuf_4
X_4349_ _4310_/A _4321_/A _4321_/B _4348_/Y vssd1 vssd1 vccd1 vccd1 _4494_/A sky130_fd_sc_hd__a31o_1
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6019_ _6020_/C _6137_/B _6020_/A _6110_/A vssd1 vssd1 vccd1 vccd1 _6021_/A sky130_fd_sc_hd__a22oi_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3720_ _3720_/A _3720_/B _3720_/C _3720_/D vssd1 vssd1 vccd1 vccd1 _3723_/A sky130_fd_sc_hd__nand4_1
X_3651_ _4407_/A vssd1 vssd1 vccd1 vccd1 _4068_/A sky130_fd_sc_hd__buf_2
X_3582_ _3607_/B _3607_/C _3582_/C vssd1 vssd1 vccd1 vccd1 _3586_/C sky130_fd_sc_hd__nand3_4
X_5321_ _5328_/A _5321_/B _5321_/C vssd1 vssd1 vccd1 vccd1 _5321_/X sky130_fd_sc_hd__and3_1
X_5252_ _5263_/A _5263_/B _5248_/Y vssd1 vssd1 vccd1 vccd1 _5252_/X sky130_fd_sc_hd__a21o_1
X_5183_ _5182_/A _5182_/B _5182_/C vssd1 vssd1 vccd1 vccd1 _5184_/C sky130_fd_sc_hd__a21o_1
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4203_ input4/X vssd1 vssd1 vccd1 vccd1 _4708_/C sky130_fd_sc_hd__buf_2
X_4134_ _3873_/Y _3872_/Y _4220_/A _4135_/B _4115_/Y vssd1 vssd1 vccd1 vccd1 _4134_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4065_ _4065_/A vssd1 vssd1 vccd1 vccd1 _5284_/C sky130_fd_sc_hd__buf_4
XFILLER_83_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4967_ _4957_/X _4955_/Y _4959_/Y _4954_/Y _4948_/Y vssd1 vssd1 vccd1 vccd1 _4968_/C
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3918_ _3918_/A _3918_/B _3918_/C vssd1 vssd1 vccd1 vccd1 _3918_/X sky130_fd_sc_hd__and3_1
X_4898_ _4898_/A _5113_/A _5113_/B vssd1 vssd1 vccd1 vccd1 _4981_/C sky130_fd_sc_hd__nand3_2
X_3849_ _3999_/A _3845_/A _3729_/C _3848_/Y vssd1 vssd1 vccd1 vccd1 _3849_/Y sky130_fd_sc_hd__o2bb2ai_2
X_5519_ _5519_/A _5519_/B _5519_/C vssd1 vssd1 vccd1 vccd1 _5519_/X sky130_fd_sc_hd__and3_1
XFILLER_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5870_ _5912_/A _5869_/Y _5859_/Y vssd1 vssd1 vccd1 vccd1 _5870_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_80_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4821_ _4822_/B _4822_/C _4822_/A vssd1 vssd1 vccd1 vccd1 _4824_/A sky130_fd_sc_hd__a21o_1
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4752_ _4752_/A vssd1 vssd1 vccd1 vccd1 _4890_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4683_ _4683_/A _4683_/B _4683_/C vssd1 vssd1 vccd1 vccd1 _4842_/D sky130_fd_sc_hd__nand3_1
X_3703_ _3703_/A _3703_/B vssd1 vssd1 vccd1 vccd1 _3703_/Y sky130_fd_sc_hd__nand2_1
X_3634_ _3634_/A vssd1 vssd1 vccd1 vccd1 _3634_/X sky130_fd_sc_hd__clkbuf_8
X_3565_ _3565_/A _3565_/B vssd1 vssd1 vccd1 vccd1 _3565_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5304_ _5304_/A _5304_/B vssd1 vssd1 vccd1 vccd1 _5307_/A sky130_fd_sc_hd__nand2_1
X_6284_ _6259_/X _6281_/Y _6283_/X vssd1 vssd1 vccd1 vccd1 _6286_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3496_ _4901_/A vssd1 vssd1 vccd1 vccd1 _5655_/A sky130_fd_sc_hd__clkbuf_4
X_5235_ _5060_/Y _5081_/B _5234_/Y vssd1 vssd1 vccd1 vccd1 _5236_/B sky130_fd_sc_hd__a21oi_4
X_5166_ _5178_/A _5178_/B _5177_/A vssd1 vssd1 vccd1 vccd1 _5171_/D sky130_fd_sc_hd__nand3_1
XFILLER_68_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5097_ _5202_/A vssd1 vssd1 vccd1 vccd1 _5278_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4117_ _4211_/B vssd1 vssd1 vccd1 vccd1 _4127_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4048_ _4681_/A _4048_/B _4048_/C vssd1 vssd1 vccd1 vccd1 _4048_/Y sky130_fd_sc_hd__nand3_1
X_5999_ _6090_/C _5999_/B vssd1 vssd1 vccd1 vccd1 _5999_/X sky130_fd_sc_hd__or2_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3350_ _4547_/A vssd1 vssd1 vccd1 vccd1 _3350_/Y sky130_fd_sc_hd__clkinv_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5020_/A _5020_/B vssd1 vssd1 vccd1 vccd1 _5020_/Y sky130_fd_sc_hd__nand2_2
XFILLER_2_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3281_ _3345_/B _3287_/A _4747_/A _3280_/X vssd1 vssd1 vccd1 vccd1 _3295_/A sky130_fd_sc_hd__o2bb2ai_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5922_ _5927_/A _6137_/C _6132_/C _5927_/C vssd1 vssd1 vccd1 vccd1 _6025_/B sky130_fd_sc_hd__nand4_1
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5853_ _5850_/X _5852_/X _5848_/Y _5840_/Y vssd1 vssd1 vccd1 vccd1 _5853_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5784_ _5884_/A _5766_/C _5766_/B vssd1 vssd1 vccd1 vccd1 _5883_/A sky130_fd_sc_hd__a21bo_1
X_4804_ _4793_/X _4798_/Y _4803_/Y vssd1 vssd1 vccd1 vccd1 _4814_/A sky130_fd_sc_hd__o21ai_1
X_4735_ _5065_/B vssd1 vssd1 vccd1 vccd1 _6171_/A sky130_fd_sc_hd__clkinv_4
X_4666_ _4678_/A vssd1 vssd1 vccd1 vccd1 _4680_/C sky130_fd_sc_hd__buf_2
X_3617_ _3617_/A vssd1 vssd1 vccd1 vccd1 _3806_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4597_ _4597_/A _4597_/B vssd1 vssd1 vccd1 vccd1 _4598_/A sky130_fd_sc_hd__nand2_2
X_3548_ _3461_/Y _3525_/Y _3458_/Y vssd1 vssd1 vccd1 vccd1 _3565_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6267_ _6277_/A _6275_/B vssd1 vssd1 vccd1 vccd1 _6267_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3479_ _3479_/A _3486_/A _3486_/B vssd1 vssd1 vccd1 vccd1 _3479_/Y sky130_fd_sc_hd__nand3_1
XFILLER_88_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5218_ _5218_/A _5218_/B _5218_/C vssd1 vssd1 vccd1 vccd1 _5271_/A sky130_fd_sc_hd__nand3_1
X_6198_ _6198_/A _6173_/C vssd1 vssd1 vccd1 vccd1 _6213_/A sky130_fd_sc_hd__or2b_1
X_5149_ _5149_/A vssd1 vssd1 vccd1 vccd1 _5163_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4520_ _4520_/A _4520_/B vssd1 vssd1 vccd1 vccd1 _4520_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4451_ _3474_/A _5453_/A _4476_/A vssd1 vssd1 vccd1 vccd1 _4451_/X sky130_fd_sc_hd__o21a_1
X_3402_ _3514_/A _5833_/A vssd1 vssd1 vccd1 vccd1 _3402_/Y sky130_fd_sc_hd__nand2_1
X_6121_ _6108_/A _6108_/B _6108_/C _6159_/B vssd1 vssd1 vccd1 vccd1 _6121_/Y sky130_fd_sc_hd__a31oi_2
X_4382_ _4110_/Y _4105_/B _4109_/Y vssd1 vssd1 vccd1 vccd1 _4382_/X sky130_fd_sc_hd__a21o_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _5373_/A vssd1 vssd1 vccd1 vccd1 _5596_/B sky130_fd_sc_hd__clkbuf_4
X_6052_ _5933_/B _5987_/Y _6054_/A vssd1 vssd1 vccd1 vccd1 _6058_/B sky130_fd_sc_hd__a21o_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _4593_/A vssd1 vssd1 vccd1 vccd1 _5263_/C sky130_fd_sc_hd__buf_4
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _4723_/X _4809_/B _4986_/X _4991_/Y vssd1 vssd1 vccd1 vccd1 _5005_/B sky130_fd_sc_hd__o22ai_2
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _3772_/A vssd1 vssd1 vccd1 vccd1 _5066_/A sky130_fd_sc_hd__buf_2
XFILLER_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5905_ _5905_/A _5905_/B _6065_/D _6127_/D vssd1 vssd1 vccd1 vccd1 _5998_/A sky130_fd_sc_hd__nand4_4
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5836_ _5905_/B _6127_/C vssd1 vssd1 vccd1 vccd1 _6096_/A sky130_fd_sc_hd__nand2_1
X_5767_ _5527_/A _5634_/C _5634_/D vssd1 vssd1 vccd1 vccd1 _5768_/C sky130_fd_sc_hd__a21boi_1
X_5698_ _5919_/A _5794_/B _5931_/A _5794_/C vssd1 vssd1 vccd1 vccd1 _5698_/Y sky130_fd_sc_hd__nand4_2
X_4718_ _4722_/A _4988_/A _4722_/B vssd1 vssd1 vccd1 vccd1 _4988_/B sky130_fd_sc_hd__nand3_1
X_4649_ _4643_/A _4643_/B _4631_/A _4631_/B vssd1 vssd1 vccd1 vccd1 _4649_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_76_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3951_ _4186_/B vssd1 vssd1 vccd1 vccd1 _6165_/B sky130_fd_sc_hd__buf_2
XFILLER_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3882_ _3980_/B _3882_/B _3882_/C vssd1 vssd1 vccd1 vccd1 _3938_/B sky130_fd_sc_hd__and3_1
XFILLER_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5621_ _5619_/Y _5620_/X _5625_/A _5625_/B vssd1 vssd1 vccd1 vccd1 _5622_/C sky130_fd_sc_hd__o211ai_2
X_5552_ _5034_/B _5453_/B _5538_/X _5540_/X _5542_/Y vssd1 vssd1 vccd1 vccd1 _5555_/B
+ sky130_fd_sc_hd__o221ai_4
X_4503_ _4323_/B _4323_/C _4323_/A vssd1 vssd1 vccd1 vccd1 _4503_/Y sky130_fd_sc_hd__a21oi_1
X_5483_ _5483_/A _5483_/B _5483_/C vssd1 vssd1 vccd1 vccd1 _5502_/A sky130_fd_sc_hd__nand3_2
XFILLER_6_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4434_ _4600_/A _4600_/B _4600_/C vssd1 vssd1 vccd1 vccd1 _4601_/A sky130_fd_sc_hd__a21o_1
X_4365_ _4365_/A _4365_/B vssd1 vssd1 vccd1 vccd1 _4365_/Y sky130_fd_sc_hd__nand2_2
X_6104_ _6104_/A _6104_/B _6104_/C vssd1 vssd1 vccd1 vccd1 _6108_/B sky130_fd_sc_hd__nand3_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ _3315_/A _3598_/A _3315_/C vssd1 vssd1 vccd1 vccd1 _3317_/B sky130_fd_sc_hd__a21oi_1
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6035_ _5999_/X _6035_/B _6035_/C vssd1 vssd1 vccd1 vccd1 _6041_/A sky130_fd_sc_hd__nand3b_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _4296_/A vssd1 vssd1 vccd1 vccd1 _4308_/A sky130_fd_sc_hd__clkbuf_2
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _3170_/A _3170_/B _3202_/B _3245_/B _6297_/A vssd1 vssd1 vccd1 vccd1 _3598_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3178_ _4708_/A vssd1 vssd1 vccd1 vccd1 _4941_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5819_ _5728_/A _5733_/Y _5726_/Y vssd1 vssd1 vccd1 vccd1 _5865_/C sky130_fd_sc_hd__a21oi_2
XFILLER_22_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4150_ _4150_/A _4150_/B _4150_/C vssd1 vssd1 vccd1 vccd1 _4151_/A sky130_fd_sc_hd__nand3_1
X_4081_ _4064_/X _4079_/Y _3223_/B _4080_/X _4071_/Y vssd1 vssd1 vccd1 vccd1 _4284_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4983_ _4980_/Y _4982_/Y _4972_/Y vssd1 vssd1 vccd1 vccd1 _4985_/A sky130_fd_sc_hd__o21ai_1
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3934_ _3934_/A _3934_/B vssd1 vssd1 vccd1 vccd1 _3934_/Y sky130_fd_sc_hd__nand2_2
X_3865_ _3867_/A _5211_/A vssd1 vssd1 vccd1 vccd1 _4103_/A sky130_fd_sc_hd__nand2_4
X_5604_ _5604_/A _5604_/B _5661_/A vssd1 vssd1 vccd1 vccd1 _5604_/X sky130_fd_sc_hd__and3_1
X_3796_ _3791_/A _3791_/B _3795_/Y vssd1 vssd1 vccd1 vccd1 _3799_/B sky130_fd_sc_hd__a21o_1
X_5535_ _5449_/A _5436_/B _5434_/D _5436_/A vssd1 vssd1 vccd1 vccd1 _5535_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5466_ _5465_/C _4829_/A _5640_/A _5465_/A vssd1 vssd1 vccd1 vccd1 _5468_/B sky130_fd_sc_hd__a22o_1
X_4417_ _4417_/A vssd1 vssd1 vccd1 vccd1 _4417_/X sky130_fd_sc_hd__buf_4
X_5397_ _5397_/A _5397_/B vssd1 vssd1 vccd1 vccd1 _5403_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4348_ _4309_/B _4309_/C _4309_/A vssd1 vssd1 vccd1 vccd1 _4348_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4279_ _4279_/A _4279_/B _4279_/C vssd1 vssd1 vccd1 vccd1 _4294_/B sky130_fd_sc_hd__nand3_2
X_6018_ _6079_/A _6077_/A _6076_/A _6076_/B vssd1 vssd1 vccd1 vccd1 _6110_/A sky130_fd_sc_hd__nand4_4
XFILLER_27_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3650_ _5048_/A _5123_/A vssd1 vssd1 vccd1 vccd1 _3650_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3581_ _3607_/B _3607_/C _3582_/C vssd1 vssd1 vccd1 vccd1 _3586_/B sky130_fd_sc_hd__a21o_2
X_5320_ _5321_/B _5321_/C _5328_/A vssd1 vssd1 vccd1 vccd1 _5320_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5251_ _5251_/A _5373_/A _5575_/B _5372_/C vssd1 vssd1 vccd1 vccd1 _5263_/B sky130_fd_sc_hd__nand4_4
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4202_ _4202_/A vssd1 vssd1 vccd1 vccd1 _4516_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5182_ _5182_/A _5182_/B _5182_/C vssd1 vssd1 vccd1 vccd1 _5184_/B sky130_fd_sc_hd__nand3_2
XFILLER_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4133_ _4133_/A _4133_/B vssd1 vssd1 vccd1 vccd1 _4137_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4064_ _4064_/A vssd1 vssd1 vccd1 vccd1 _4064_/X sky130_fd_sc_hd__buf_2
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4966_ _4942_/Y _4943_/X _4938_/Y _4965_/X vssd1 vssd1 vccd1 vccd1 _4968_/B sky130_fd_sc_hd__o22ai_1
XFILLER_11_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3917_ _3915_/Y _3898_/X _4890_/C _3714_/D vssd1 vssd1 vccd1 vccd1 _3917_/X sky130_fd_sc_hd__o211a_1
X_4897_ _4879_/Y _4882_/X _4865_/Y _4871_/X vssd1 vssd1 vccd1 vccd1 _5113_/B sky130_fd_sc_hd__o211ai_2
X_3848_ _3848_/A vssd1 vssd1 vccd1 vccd1 _3848_/Y sky130_fd_sc_hd__inv_2
X_3779_ _3685_/A _3685_/C _3708_/Y _3707_/X vssd1 vssd1 vccd1 vccd1 _3819_/B sky130_fd_sc_hd__o2bb2ai_2
X_5518_ _5518_/A _5518_/B _5518_/C vssd1 vssd1 vccd1 vccd1 _5980_/B sky130_fd_sc_hd__nor3_4
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5449_ _5449_/A vssd1 vssd1 vccd1 vccd1 _5712_/A sky130_fd_sc_hd__buf_2
XFILLER_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4820_ _4559_/A _4559_/B _4559_/C _4659_/B vssd1 vssd1 vccd1 vccd1 _4822_/A sky130_fd_sc_hd__a31o_2
XFILLER_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4751_ _4751_/A _4751_/B vssd1 vssd1 vccd1 vccd1 _4752_/A sky130_fd_sc_hd__nand2_1
X_4682_ _4681_/X _4508_/Y _4516_/B vssd1 vssd1 vccd1 vccd1 _4683_/C sky130_fd_sc_hd__o21ai_1
X_3702_ _3702_/A _3702_/B vssd1 vssd1 vccd1 vccd1 _3702_/Y sky130_fd_sc_hd__nand2_1
X_3633_ _3633_/A vssd1 vssd1 vccd1 vccd1 _3634_/A sky130_fd_sc_hd__clkbuf_4
X_3564_ _3564_/A _3564_/B _3564_/C vssd1 vssd1 vccd1 vccd1 _3564_/X sky130_fd_sc_hd__and3_1
XFILLER_88_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6283_ _6283_/A _6283_/B _6283_/C vssd1 vssd1 vccd1 vccd1 _6283_/X sky130_fd_sc_hd__and3_1
X_5303_ _5303_/A _5303_/B vssd1 vssd1 vccd1 vccd1 _5304_/B sky130_fd_sc_hd__nor2_1
X_3495_ _4193_/A _3960_/B _5580_/A _5404_/B vssd1 vssd1 vccd1 vccd1 _3508_/D sky130_fd_sc_hd__nand4_4
XFILLER_88_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5234_ _5240_/A _5378_/B _5240_/D _4067_/A vssd1 vssd1 vccd1 vccd1 _5234_/Y sky130_fd_sc_hd__a22oi_2
X_5165_ _5151_/Y _5153_/X _5325_/A _5157_/B vssd1 vssd1 vccd1 vccd1 _5177_/A sky130_fd_sc_hd__o211ai_2
X_4116_ _3873_/Y _3872_/Y _4115_/Y vssd1 vssd1 vccd1 vccd1 _4211_/B sky130_fd_sc_hd__a21oi_1
X_5096_ _5096_/A _5096_/B _5096_/C vssd1 vssd1 vccd1 vccd1 _5202_/A sky130_fd_sc_hd__nand3_1
XFILLER_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4047_ _4047_/A vssd1 vssd1 vccd1 vccd1 _4681_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _5998_/A _5998_/B _5998_/C vssd1 vssd1 vccd1 vccd1 _5999_/B sky130_fd_sc_hd__and3_1
XFILLER_24_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4949_ _4942_/Y _4943_/X _4948_/Y vssd1 vssd1 vccd1 vccd1 _4949_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_24_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3280_ _3280_/A vssd1 vssd1 vccd1 vccd1 _3280_/X sky130_fd_sc_hd__buf_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5921_ _6132_/C _6137_/C _5927_/C _5927_/A vssd1 vssd1 vccd1 vccd1 _6025_/A sky130_fd_sc_hd__a22o_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5852_ _5852_/A _6134_/C _5852_/C vssd1 vssd1 vccd1 vccd1 _5852_/X sky130_fd_sc_hd__and3_1
X_5783_ _5712_/A _5933_/C _5506_/X _6255_/A _5729_/B vssd1 vssd1 vccd1 vccd1 _5892_/A
+ sky130_fd_sc_hd__a41o_2
XFILLER_21_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4803_ _4803_/A _4803_/B _4803_/C vssd1 vssd1 vccd1 vccd1 _4803_/Y sky130_fd_sc_hd__nand3_1
X_4734_ _5048_/A _4734_/B _5068_/D _5245_/B vssd1 vssd1 vccd1 vccd1 _4746_/B sky130_fd_sc_hd__nand4_4
X_4665_ _4665_/A _4665_/B _4665_/C vssd1 vssd1 vccd1 vccd1 _4678_/A sky130_fd_sc_hd__nand3_1
X_4596_ _4473_/X _4592_/B _4880_/A _4080_/X _4595_/X vssd1 vssd1 vccd1 vccd1 _4597_/B
+ sky130_fd_sc_hd__o2111ai_1
X_3616_ _3616_/A _3616_/B vssd1 vssd1 vccd1 vccd1 _3617_/A sky130_fd_sc_hd__nand2_1
X_3547_ _3564_/A _3564_/B _5382_/C _5347_/A vssd1 vssd1 vccd1 vccd1 _3549_/B sky130_fd_sc_hd__nand4_1
XFILLER_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6266_ _6266_/A _6266_/B _6266_/C vssd1 vssd1 vccd1 vccd1 _6275_/B sky130_fd_sc_hd__and3_1
X_3478_ _3478_/A _3478_/B _3478_/C vssd1 vssd1 vccd1 vccd1 _3486_/B sky130_fd_sc_hd__nand3_2
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6197_ _6197_/A _6197_/B vssd1 vssd1 vccd1 vccd1 _6197_/X sky130_fd_sc_hd__xor2_4
X_5217_ _5070_/A _5204_/Y _5080_/B vssd1 vssd1 vccd1 vccd1 _5218_/C sky130_fd_sc_hd__o21ai_4
XFILLER_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5148_ _5099_/Y _4912_/Y _5146_/X _5366_/B vssd1 vssd1 vccd1 vccd1 _5149_/A sky130_fd_sc_hd__o211ai_2
X_5079_ _5211_/B vssd1 vssd1 vccd1 vccd1 _5794_/C sky130_fd_sc_hd__buf_2
XFILLER_28_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4450_ _4257_/Y _4592_/A _4449_/Y _4254_/B vssd1 vssd1 vccd1 vccd1 _4476_/A sky130_fd_sc_hd__o2bb2ai_1
X_4381_ _3448_/X _3512_/X _4103_/B _4411_/A _4422_/A vssd1 vssd1 vccd1 vccd1 _4381_/Y
+ sky130_fd_sc_hd__o221ai_4
X_3401_ _3620_/C vssd1 vssd1 vccd1 vccd1 _5833_/A sky130_fd_sc_hd__buf_4
X_6120_ _6017_/A _6017_/B _6110_/B vssd1 vssd1 vccd1 vccd1 _6159_/B sky130_fd_sc_hd__o21a_1
X_3332_ _4873_/A vssd1 vssd1 vccd1 vccd1 _5373_/A sky130_fd_sc_hd__clkbuf_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _6051_/A _6051_/B vssd1 vssd1 vccd1 vccd1 _6054_/A sky130_fd_sc_hd__nand2_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3322_/A vssd1 vssd1 vccd1 vccd1 _4593_/A sky130_fd_sc_hd__buf_2
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _4822_/A _4822_/C _4822_/B vssd1 vssd1 vccd1 vccd1 _5005_/A sky130_fd_sc_hd__a21boi_4
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3194_ input9/X vssd1 vssd1 vccd1 vccd1 _3772_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5904_ _5905_/B _6127_/C _6127_/D _5850_/A vssd1 vssd1 vccd1 vccd1 _5907_/A sky130_fd_sc_hd__a22o_1
X_5835_ _5846_/A _5846_/B _5847_/B vssd1 vssd1 vccd1 vccd1 _5840_/A sky130_fd_sc_hd__a21o_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5766_ _5884_/A _5766_/B _5766_/C vssd1 vssd1 vccd1 vccd1 _5768_/B sky130_fd_sc_hd__nand3_1
X_5697_ _5697_/A _5697_/B vssd1 vssd1 vccd1 vccd1 _5799_/A sky130_fd_sc_hd__nand2_1
X_4717_ _4711_/B _4715_/X _4716_/Y vssd1 vssd1 vccd1 vccd1 _4722_/B sky130_fd_sc_hd__o21ai_4
X_4648_ _4648_/A _4648_/B vssd1 vssd1 vccd1 vccd1 _4652_/B sky130_fd_sc_hd__nand2_2
XFILLER_30_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4579_ _4734_/B _4877_/D _5068_/D _4432_/A vssd1 vssd1 vccd1 vccd1 _4579_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6249_ _6225_/Y _6226_/X _6275_/C vssd1 vssd1 vccd1 vccd1 _6251_/A sky130_fd_sc_hd__a21oi_1
XFILLER_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3950_ _5704_/B vssd1 vssd1 vccd1 vccd1 _4186_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_16_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3881_ _3980_/B _3882_/B _3882_/C vssd1 vssd1 vccd1 vccd1 _3938_/A sky130_fd_sc_hd__a21oi_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5620_ _5612_/X _5613_/Y _5614_/Y _5611_/A _5611_/B vssd1 vssd1 vccd1 vccd1 _5620_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_31_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5551_ _5291_/X _5542_/A _5546_/Y _5547_/Y vssd1 vssd1 vccd1 vccd1 _5555_/A sky130_fd_sc_hd__o22a_1
X_4502_ _4502_/A _4502_/B _4502_/C vssd1 vssd1 vccd1 vccd1 _4506_/B sky130_fd_sc_hd__nand3_1
X_5482_ _5634_/B _5480_/Y _5477_/A _5492_/B vssd1 vssd1 vccd1 vccd1 _5483_/C sky130_fd_sc_hd__o211ai_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4433_ _4868_/A _5029_/B vssd1 vssd1 vccd1 vccd1 _4600_/C sky130_fd_sc_hd__and2_1
X_4364_ _4530_/A _4530_/C vssd1 vssd1 vccd1 vccd1 _4365_/B sky130_fd_sc_hd__nand2_2
X_6103_ _6104_/B _6104_/C _6104_/A vssd1 vssd1 vccd1 vccd1 _6108_/A sky130_fd_sc_hd__a21o_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4295_ _4295_/A _4295_/B _4295_/C vssd1 vssd1 vccd1 vccd1 _4296_/A sky130_fd_sc_hd__nand3_1
X_3315_ _3315_/A _3598_/A _3315_/C vssd1 vssd1 vccd1 vccd1 _3317_/A sky130_fd_sc_hd__and3_1
X_6034_ _6037_/A _6034_/B vssd1 vssd1 vccd1 vccd1 _6035_/C sky130_fd_sc_hd__nand2_1
XFILLER_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _3246_/A _3246_/B vssd1 vssd1 vccd1 vccd1 _3315_/A sky130_fd_sc_hd__or2_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3177_ _4019_/A vssd1 vssd1 vccd1 vccd1 _4708_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5818_ _5818_/A _5818_/B _5818_/C vssd1 vssd1 vccd1 vccd1 _5865_/B sky130_fd_sc_hd__nand3_2
XFILLER_10_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5749_ _5734_/Y _5738_/Y _5739_/X vssd1 vssd1 vccd1 vccd1 _5749_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_1_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4080_ _4777_/D vssd1 vssd1 vccd1 vccd1 _4080_/X sky130_fd_sc_hd__buf_4
XFILLER_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4982_ _4765_/B _4924_/Y _4925_/Y _4981_/Y vssd1 vssd1 vccd1 vccd1 _4982_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3933_ _3626_/X _3803_/X _3793_/Y _3799_/Y _3806_/A vssd1 vssd1 vccd1 vccd1 _3934_/B
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_51_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3864_ _3676_/B _3902_/A _3770_/Y _3768_/Y vssd1 vssd1 vccd1 vccd1 _3878_/C sky130_fd_sc_hd__o22ai_4
X_5603_ _5603_/A _6236_/B _5603_/C vssd1 vssd1 vccd1 vccd1 _5603_/X sky130_fd_sc_hd__or3_1
X_3795_ _3803_/A _3795_/B vssd1 vssd1 vccd1 vccd1 _3795_/Y sky130_fd_sc_hd__nand2_1
X_5534_ _5534_/A _5809_/B vssd1 vssd1 vccd1 vccd1 _5534_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5465_ _5465_/A _5933_/D _5465_/C _5640_/A vssd1 vssd1 vccd1 vccd1 _5640_/B sky130_fd_sc_hd__nand4_2
X_4416_ _4406_/Y _4408_/Y _4251_/Y vssd1 vssd1 vccd1 vccd1 _4416_/Y sky130_fd_sc_hd__o21ai_1
X_5396_ _5236_/A _5236_/B _5612_/A _5612_/B _5395_/Y vssd1 vssd1 vccd1 vccd1 _5614_/A
+ sky130_fd_sc_hd__o2111ai_4
X_4347_ _4832_/C _6255_/A vssd1 vssd1 vccd1 vccd1 _4681_/B sky130_fd_sc_hd__nand2_4
X_4278_ _4059_/Y _4063_/Y _4073_/Y vssd1 vssd1 vccd1 vccd1 _4279_/C sky130_fd_sc_hd__o21ai_1
XFILLER_74_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6017_ _6017_/A _6017_/B vssd1 vssd1 vccd1 vccd1 _6020_/A sky130_fd_sc_hd__nand2_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3229_ _3229_/A _3229_/B _4827_/A _3229_/D vssd1 vssd1 vccd1 vccd1 _3230_/B sky130_fd_sc_hd__nand4_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3580_ _3402_/Y _3498_/A _3407_/X _3410_/B vssd1 vssd1 vccd1 vccd1 _3582_/C sky130_fd_sc_hd__o211a_2
XFILLER_42_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5250_ _5250_/A _5250_/B vssd1 vssd1 vccd1 vccd1 _5263_/A sky130_fd_sc_hd__nand2_4
X_4201_ _4201_/A _5805_/B _4201_/C vssd1 vssd1 vccd1 vccd1 _4202_/A sky130_fd_sc_hd__and3_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5181_ _3280_/X _6235_/A _4955_/Y _4943_/B vssd1 vssd1 vccd1 vccd1 _5182_/C sky130_fd_sc_hd__o31a_1
XFILLER_95_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4132_ _4126_/Y _4127_/X _4130_/Y _4131_/Y vssd1 vssd1 vccd1 vccd1 _4137_/A sky130_fd_sc_hd__o22ai_4
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4063_ _5053_/A _5206_/A _4884_/B _5048_/A vssd1 vssd1 vccd1 vccd1 _4063_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_95_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4965_ _4703_/X _4944_/X _4946_/Y _4947_/X vssd1 vssd1 vccd1 vccd1 _4965_/X sky130_fd_sc_hd__o22a_2
X_3916_ _5064_/A vssd1 vssd1 vccd1 vccd1 _4890_/C sky130_fd_sc_hd__buf_4
XFILLER_32_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4896_ _4865_/Y _4871_/X _4885_/X _4886_/Y vssd1 vssd1 vccd1 vccd1 _5113_/A sky130_fd_sc_hd__o2bb2ai_1
X_3847_ _3847_/A _3847_/B _3847_/C vssd1 vssd1 vccd1 vccd1 _3999_/A sky130_fd_sc_hd__nand3_2
X_3778_ _3778_/A _3809_/B vssd1 vssd1 vccd1 vccd1 _3819_/A sky130_fd_sc_hd__nand2_1
X_5517_ _5517_/A _5520_/A _5520_/B _5517_/D vssd1 vssd1 vccd1 vccd1 _5518_/C sky130_fd_sc_hd__nand4_4
X_5448_ _5448_/A _5448_/B vssd1 vssd1 vccd1 vccd1 _5542_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5379_ _5379_/A vssd1 vssd1 vccd1 vccd1 _5598_/A sky130_fd_sc_hd__buf_2
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4750_ _4877_/A _4873_/B vssd1 vssd1 vccd1 vccd1 _4751_/B sky130_fd_sc_hd__nand2_1
X_4681_ _4681_/A _4681_/B vssd1 vssd1 vccd1 vccd1 _4681_/X sky130_fd_sc_hd__or2_1
X_3701_ _3688_/X _3689_/Y _3687_/A _3690_/Y _3700_/Y vssd1 vssd1 vccd1 vccd1 _3705_/B
+ sky130_fd_sc_hd__o221ai_2
X_3632_ _3632_/A _3632_/B _3632_/C vssd1 vssd1 vccd1 vccd1 _3691_/A sky130_fd_sc_hd__nand3_2
X_5302_ _5511_/A _5302_/B _5302_/C _5514_/A vssd1 vssd1 vccd1 vccd1 _5303_/B sky130_fd_sc_hd__and4_2
X_3563_ _3465_/Y _3446_/A _3462_/Y _3459_/Y vssd1 vssd1 vccd1 vccd1 _3567_/B sky130_fd_sc_hd__o2bb2ai_1
X_6282_ _5967_/X _6255_/C _6258_/A _6258_/B vssd1 vssd1 vccd1 vccd1 _6283_/A sky130_fd_sc_hd__a22o_1
X_3494_ _5026_/B vssd1 vssd1 vccd1 vccd1 _5404_/B sky130_fd_sc_hd__buf_4
X_5233_ _5258_/A _5229_/Y _5232_/Y vssd1 vssd1 vccd1 vccd1 _5236_/A sky130_fd_sc_hd__o21a_2
X_5164_ _5325_/A _5157_/B _5161_/X _5163_/X vssd1 vssd1 vccd1 vccd1 _5178_/B sky130_fd_sc_hd__o2bb2ai_1
X_4115_ _5302_/C _5663_/A _5663_/B _5134_/A vssd1 vssd1 vccd1 vccd1 _4115_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5095_ _5095_/A _5095_/B _5257_/A _5257_/B vssd1 vssd1 vccd1 vccd1 _5096_/C sky130_fd_sc_hd__nand4_1
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4046_ _4362_/C _6016_/A vssd1 vssd1 vccd1 vccd1 _4047_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5997_ _5998_/A _5998_/B _5998_/C vssd1 vssd1 vccd1 vccd1 _6090_/C sky130_fd_sc_hd__a21oi_2
XFILLER_33_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4948_ _4703_/X _4944_/X _4946_/Y _4947_/X vssd1 vssd1 vccd1 vccd1 _4948_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_20_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4879_ _5678_/B _5407_/C _4885_/B _4885_/C vssd1 vssd1 vccd1 vccd1 _4879_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5920_ _5920_/A _5920_/B vssd1 vssd1 vccd1 vccd1 _5927_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5851_ _6010_/B vssd1 vssd1 vccd1 vccd1 _6134_/C sky130_fd_sc_hd__clkbuf_2
X_5782_ _5782_/A _5782_/B vssd1 vssd1 vccd1 vccd1 _5891_/A sky130_fd_sc_hd__nand2_1
X_4802_ _4802_/A _4802_/B vssd1 vssd1 vccd1 vccd1 _4803_/C sky130_fd_sc_hd__nand2_1
X_4733_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5245_/B sky130_fd_sc_hd__buf_2
X_4664_ _4653_/A _4663_/B _4669_/A vssd1 vssd1 vccd1 vccd1 _4665_/C sky130_fd_sc_hd__a21o_1
X_3615_ _4026_/A _5026_/A vssd1 vssd1 vccd1 vccd1 _3616_/B sky130_fd_sc_hd__nand2_1
X_4595_ _5065_/A _5206_/A _5539_/B _5066_/A vssd1 vssd1 vccd1 vccd1 _4595_/X sky130_fd_sc_hd__a22o_1
X_3546_ _4945_/A vssd1 vssd1 vccd1 vccd1 _5347_/A sky130_fd_sc_hd__clkbuf_4
X_6265_ _6266_/A _6266_/C _6266_/B vssd1 vssd1 vccd1 vccd1 _6277_/A sky130_fd_sc_hd__a21oi_1
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5216_ _5025_/B _5403_/A _4110_/B _5704_/A _5208_/Y vssd1 vssd1 vccd1 vccd1 _5218_/B
+ sky130_fd_sc_hd__o2111ai_4
X_3477_ _3477_/A _3477_/B vssd1 vssd1 vccd1 vccd1 _3478_/C sky130_fd_sc_hd__nand2_1
X_6196_ _5982_/B _6193_/Y _6195_/Y vssd1 vssd1 vccd1 vccd1 _6197_/B sky130_fd_sc_hd__a21oi_4
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5147_ _5140_/Y _5141_/X _5126_/Y _5366_/A vssd1 vssd1 vccd1 vccd1 _5366_/B sky130_fd_sc_hd__o211ai_4
XFILLER_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5078_ _5594_/A _5925_/B _5080_/A _5070_/C vssd1 vssd1 vccd1 vccd1 _5078_/Y sky130_fd_sc_hd__a22oi_2
X_4029_ _4176_/A _5553_/B vssd1 vssd1 vccd1 vccd1 _4029_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4380_ _4693_/A _5029_/A vssd1 vssd1 vccd1 vccd1 _4411_/A sky130_fd_sc_hd__nand2_2
X_3400_ _5397_/A vssd1 vssd1 vccd1 vccd1 _3620_/C sky130_fd_sc_hd__clkbuf_2
X_3331_ _3897_/A vssd1 vssd1 vccd1 vccd1 _4873_/A sky130_fd_sc_hd__clkbuf_4
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _5960_/X _5964_/Y _6048_/A _6048_/B vssd1 vssd1 vccd1 vccd1 _6051_/B sky130_fd_sc_hd__o211ai_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3265_/D _3265_/A _3186_/A _5390_/A vssd1 vssd1 vccd1 vccd1 _3306_/A sky130_fd_sc_hd__o2bb2ai_2
X_5001_ _5020_/A _5020_/B _5001_/C vssd1 vssd1 vccd1 vccd1 _5001_/Y sky130_fd_sc_hd__nand3_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ _3242_/A _3242_/B _3242_/C vssd1 vssd1 vccd1 vccd1 _3199_/B sky130_fd_sc_hd__nand3_1
X_5903_ _6170_/D vssd1 vssd1 vccd1 vccd1 _6203_/C sky130_fd_sc_hd__clkbuf_2
X_5834_ _5834_/A _6001_/C vssd1 vssd1 vccd1 vccd1 _5847_/B sky130_fd_sc_hd__and2_1
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5765_ _5634_/D _5649_/X _5763_/Y _5764_/X vssd1 vssd1 vccd1 vccd1 _5781_/A sky130_fd_sc_hd__o2bb2ai_1
X_4716_ _4711_/D _4711_/B _4714_/X vssd1 vssd1 vccd1 vccd1 _4716_/Y sky130_fd_sc_hd__o21ai_1
X_5696_ _5696_/A _5701_/B vssd1 vssd1 vccd1 vccd1 _5697_/B sky130_fd_sc_hd__nand2_1
X_4647_ _4647_/A _4647_/B vssd1 vssd1 vccd1 vccd1 _4648_/B sky130_fd_sc_hd__nand2_1
XFILLER_1_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4578_ _4578_/A vssd1 vssd1 vccd1 vccd1 _5068_/D sky130_fd_sc_hd__clkbuf_4
X_3529_ _5045_/A _3758_/B vssd1 vssd1 vccd1 vccd1 _3530_/B sky130_fd_sc_hd__nand2_2
X_6248_ _6248_/A _6248_/B vssd1 vssd1 vccd1 vccd1 _6275_/C sky130_fd_sc_hd__or2_2
X_6179_ _6180_/A _6180_/C _6180_/B vssd1 vssd1 vccd1 vccd1 _6183_/A sky130_fd_sc_hd__a21oi_4
XFILLER_57_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3880_ _3468_/A _3797_/X _3879_/Y _3791_/B vssd1 vssd1 vccd1 vccd1 _3882_/C sky130_fd_sc_hd__o31a_2
X_5550_ _5550_/A _5694_/C vssd1 vssd1 vccd1 vccd1 _5550_/Y sky130_fd_sc_hd__nand2_1
X_5481_ _5418_/Y _5426_/Y _5624_/A vssd1 vssd1 vccd1 vccd1 _5492_/B sky130_fd_sc_hd__o21ai_1
X_4501_ _4502_/A _4502_/B _4502_/C vssd1 vssd1 vccd1 vccd1 _4506_/C sky130_fd_sc_hd__a21o_1
XANTENNA_0 _4287_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4432_ _4432_/A _4734_/B _4873_/B _5397_/B vssd1 vssd1 vccd1 vccd1 _4600_/B sky130_fd_sc_hd__nand4_4
X_4363_ _4363_/A _4363_/B _5792_/A _4363_/D vssd1 vssd1 vccd1 vccd1 _4363_/Y sky130_fd_sc_hd__nand4_4
X_6102_ _6024_/Y _6022_/Y _6034_/B _6030_/Y vssd1 vssd1 vccd1 vccd1 _6104_/A sky130_fd_sc_hd__a2bb2o_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ _4298_/C _4294_/B _4294_/C vssd1 vssd1 vccd1 vccd1 _4295_/C sky130_fd_sc_hd__nand3_1
X_3314_ _3598_/B vssd1 vssd1 vccd1 vccd1 _3315_/C sky130_fd_sc_hd__clkbuf_1
X_6033_ _6025_/X _5942_/A _5942_/B vssd1 vssd1 vccd1 vccd1 _6034_/B sky130_fd_sc_hd__o21ai_2
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3245_ _3245_/A _3245_/B vssd1 vssd1 vccd1 vccd1 _3245_/Y sky130_fd_sc_hd__xnor2_4
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3176_ _3210_/A vssd1 vssd1 vccd1 vccd1 _4019_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5817_ _5673_/B _5690_/X _5673_/A vssd1 vssd1 vccd1 vccd1 _5818_/C sky130_fd_sc_hd__a21boi_1
XFILLER_10_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5748_ _5748_/A _5748_/B _5748_/C vssd1 vssd1 vccd1 vccd1 _5748_/X sky130_fd_sc_hd__and3_2
X_5679_ _6124_/B vssd1 vssd1 vccd1 vccd1 _6065_/D sky130_fd_sc_hd__buf_2
XFILLER_1_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4981_ _4981_/A _4981_/B _4981_/C vssd1 vssd1 vccd1 vccd1 _4981_/Y sky130_fd_sc_hd__nand3_1
XFILLER_51_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3932_ _3793_/Y _3799_/Y _3804_/X vssd1 vssd1 vccd1 vccd1 _3934_/A sky130_fd_sc_hd__a21o_1
X_3863_ _3833_/X _3839_/B _3823_/Y vssd1 vssd1 vccd1 vccd1 _3976_/A sky130_fd_sc_hd__a21oi_2
X_5602_ _5603_/C _5229_/Y _5601_/Y _5612_/A vssd1 vssd1 vccd1 vccd1 _5686_/B sky130_fd_sc_hd__o211ai_4
X_5533_ _5531_/Y _5532_/X _4621_/C _5718_/A vssd1 vssd1 vccd1 vccd1 _5694_/A sky130_fd_sc_hd__o211ai_2
X_3794_ _3611_/X _3679_/Y _3783_/Y _3713_/Y vssd1 vssd1 vccd1 vccd1 _3799_/A sky130_fd_sc_hd__o22a_1
X_5464_ _5464_/A vssd1 vssd1 vccd1 vccd1 _5640_/A sky130_fd_sc_hd__clkbuf_2
X_5395_ _5244_/Y _5249_/Y _5252_/X _5268_/A vssd1 vssd1 vccd1 vccd1 _5395_/Y sky130_fd_sc_hd__o211ai_2
X_4415_ _3620_/C _5532_/A _4236_/B _5399_/A _4402_/Y vssd1 vssd1 vccd1 vccd1 _4415_/X
+ sky130_fd_sc_hd__a41o_1
X_4346_ _5348_/D vssd1 vssd1 vccd1 vccd1 _6255_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4277_ _4277_/A _4277_/B _4277_/C _4761_/B vssd1 vssd1 vccd1 vccd1 _4279_/B sky130_fd_sc_hd__nand4_1
X_6016_ _6016_/A _6076_/A vssd1 vssd1 vccd1 vccd1 _6017_/B sky130_fd_sc_hd__nand2_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3228_ _3639_/A _3204_/B _3229_/A _3229_/B vssd1 vssd1 vccd1 vccd1 _3230_/A sky130_fd_sc_hd__a22o_1
X_3159_ _5087_/C vssd1 vssd1 vccd1 vccd1 _3204_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_82_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4200_ _4384_/A vssd1 vssd1 vccd1 vccd1 _5805_/B sky130_fd_sc_hd__clkbuf_4
X_5180_ _5180_/A _5180_/B _5180_/C vssd1 vssd1 vccd1 vccd1 _5182_/B sky130_fd_sc_hd__nand3_4
X_4131_ _4095_/A _4095_/B _4095_/C vssd1 vssd1 vccd1 vccd1 _4131_/Y sky130_fd_sc_hd__a21oi_4
X_4062_ _4590_/B vssd1 vssd1 vccd1 vccd1 _4884_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_76_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4964_ _4950_/A _4950_/B _4951_/A vssd1 vssd1 vccd1 vccd1 _4968_/A sky130_fd_sc_hd__a21boi_1
X_3915_ _3418_/A _4619_/B _4238_/C _4454_/B vssd1 vssd1 vccd1 vccd1 _3915_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_51_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4895_ _4891_/Y _4742_/X _4768_/Y _4769_/Y vssd1 vssd1 vccd1 vccd1 _4898_/A sky130_fd_sc_hd__o2bb2ai_1
X_3846_ _3999_/B vssd1 vssd1 vccd1 vccd1 _3996_/B sky130_fd_sc_hd__buf_2
X_3777_ _3768_/Y _3771_/X _3776_/Y vssd1 vssd1 vccd1 vccd1 _3809_/B sky130_fd_sc_hd__o21ai_2
X_5516_ _5776_/A _5776_/B vssd1 vssd1 vccd1 vccd1 _5523_/A sky130_fd_sc_hd__nand2_2
X_5447_ _5442_/Y _5445_/Y _5453_/A _6236_/A vssd1 vssd1 vccd1 vccd1 _5451_/B sky130_fd_sc_hd__o2bb2ai_1
X_5378_ _5378_/A _5378_/B vssd1 vssd1 vccd1 vccd1 _5379_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4329_ _4152_/A _4170_/X _4157_/B vssd1 vssd1 vccd1 vccd1 _4334_/A sky130_fd_sc_hd__o21ai_1
XFILLER_86_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3700_ _3696_/Y _3697_/X _3719_/A _3699_/Y vssd1 vssd1 vccd1 vccd1 _3700_/Y sky130_fd_sc_hd__o211ai_1
X_4680_ _4680_/A _4680_/B _4680_/C _4680_/D vssd1 vssd1 vccd1 vccd1 _4683_/B sky130_fd_sc_hd__nand4_1
X_3631_ _3552_/A _3611_/X _3554_/Y _3555_/Y vssd1 vssd1 vccd1 vccd1 _3632_/C sky130_fd_sc_hd__a22oi_2
X_3562_ _3540_/A _3558_/B _3560_/B vssd1 vssd1 vccd1 vccd1 _3567_/A sky130_fd_sc_hd__a21o_1
X_5301_ _4422_/C _5302_/B _5514_/A _5511_/A vssd1 vssd1 vccd1 vccd1 _5303_/A sky130_fd_sc_hd__a22oi_4
X_6281_ _6283_/C _6283_/B vssd1 vssd1 vccd1 vccd1 _6281_/Y sky130_fd_sc_hd__nand2_1
X_3493_ _4906_/A vssd1 vssd1 vccd1 vccd1 _5026_/B sky130_fd_sc_hd__buf_2
X_5232_ _5232_/A _5232_/B vssd1 vssd1 vccd1 vccd1 _5232_/Y sky130_fd_sc_hd__nand2_1
X_5163_ _5336_/A _5163_/B _5163_/C vssd1 vssd1 vccd1 vccd1 _5163_/X sky130_fd_sc_hd__and3_1
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4114_ _4109_/Y _4302_/B _4112_/X _4113_/X vssd1 vssd1 vccd1 vccd1 _4211_/A sky130_fd_sc_hd__o211ai_2
XFILLER_83_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5094_ _4875_/B _5250_/A _5093_/Y vssd1 vssd1 vccd1 vccd1 _5257_/B sky130_fd_sc_hd__o21ai_1
X_4045_ _3878_/A _3878_/B _3878_/C _3980_/A vssd1 vssd1 vccd1 vccd1 _4045_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5996_ _6143_/C _5996_/B vssd1 vssd1 vccd1 vccd1 _5998_/C sky130_fd_sc_hd__or2_1
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4947_ _4928_/X _5124_/A _4945_/X _4933_/A vssd1 vssd1 vccd1 vccd1 _4947_/X sky130_fd_sc_hd__o211a_1
X_4878_ _4878_/A vssd1 vssd1 vccd1 vccd1 _4885_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3829_ _3966_/A _3829_/B _3829_/C _6165_/A vssd1 vssd1 vccd1 vccd1 _3829_/X sky130_fd_sc_hd__and4_1
XFILLER_58_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5850_ _5850_/A _5905_/B _6071_/A _6065_/C vssd1 vssd1 vccd1 vccd1 _5850_/X sky130_fd_sc_hd__and4_2
X_5781_ _5781_/A _5781_/B vssd1 vssd1 vccd1 vccd1 _5782_/B sky130_fd_sc_hd__nand2_1
XFILLER_61_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4801_ _4801_/A _4801_/B vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__nand2_1
X_4732_ _4732_/A vssd1 vssd1 vccd1 vccd1 _5059_/A sky130_fd_sc_hd__clkbuf_2
X_4663_ _4663_/A _4663_/B _4669_/A vssd1 vssd1 vccd1 vccd1 _4665_/B sky130_fd_sc_hd__nand3_1
X_3614_ _4901_/A vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__clkbuf_4
X_4594_ _4589_/Y _4592_/Y _4593_/Y vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__o21ai_1
X_3545_ _3711_/A vssd1 vssd1 vccd1 vccd1 _4945_/A sky130_fd_sc_hd__buf_2
X_6264_ _6264_/A _6264_/B vssd1 vssd1 vccd1 vccd1 _6266_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3476_ _3475_/Y _3370_/X _3344_/Y _3349_/Y vssd1 vssd1 vccd1 vccd1 _3477_/B sky130_fd_sc_hd__o2bb2ai_1
X_5215_ _5208_/Y _5209_/Y _5034_/A _4261_/Y vssd1 vssd1 vccd1 vccd1 _5218_/A sky130_fd_sc_hd__o2bb2ai_4
X_6195_ _6219_/B _6161_/B _6193_/C _6116_/X _6194_/Y vssd1 vssd1 vccd1 vccd1 _6195_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_69_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5146_ _5126_/Y _5131_/A _5138_/Y vssd1 vssd1 vccd1 vccd1 _5146_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5077_ _5211_/B vssd1 vssd1 vccd1 vccd1 _5925_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4028_ _4936_/B vssd1 vssd1 vccd1 vccd1 _5553_/B sky130_fd_sc_hd__clkbuf_4
X_5979_ _5521_/Y _5980_/C _5978_/Y vssd1 vssd1 vccd1 vccd1 _5981_/A sky130_fd_sc_hd__a21oi_4
XFILLER_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3330_ _5374_/A vssd1 vssd1 vccd1 vccd1 _5596_/A sky130_fd_sc_hd__buf_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _4723_/X _4809_/B _5021_/B _5021_/C vssd1 vssd1 vccd1 vccd1 _5001_/C sky130_fd_sc_hd__o211ai_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _4460_/A vssd1 vssd1 vccd1 vccd1 _5390_/A sky130_fd_sc_hd__buf_2
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3192_ _3242_/A _3242_/B _3242_/C vssd1 vssd1 vccd1 vccd1 _3199_/A sky130_fd_sc_hd__a21o_1
XFILLER_78_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5902_ _6003_/B vssd1 vssd1 vccd1 vccd1 _6170_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5833_ _5833_/A _5833_/B _6003_/B _6124_/B vssd1 vssd1 vccd1 vccd1 _5846_/B sky130_fd_sc_hd__nand4_2
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5764_ _5884_/A _5766_/B _5766_/C vssd1 vssd1 vccd1 vccd1 _5764_/X sky130_fd_sc_hd__and3_1
X_5695_ _5704_/A vssd1 vssd1 vccd1 vccd1 _5809_/A sky130_fd_sc_hd__buf_2
X_4715_ _3803_/B _3783_/A _5436_/B _5434_/D _4714_/X vssd1 vssd1 vccd1 vccd1 _4715_/X
+ sky130_fd_sc_hd__a41o_1
X_4646_ _4806_/A _4817_/B _4639_/Y _4645_/Y vssd1 vssd1 vccd1 vccd1 _4652_/A sky130_fd_sc_hd__a22o_1
X_4577_ _4443_/Y _4575_/Y _4600_/B _4605_/C vssd1 vssd1 vccd1 vccd1 _4577_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3528_ _3903_/A vssd1 vssd1 vccd1 vccd1 _3758_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6247_ _6247_/A _6247_/B vssd1 vssd1 vccd1 vccd1 _6248_/B sky130_fd_sc_hd__and2_1
X_3459_ _3204_/B _4422_/C _3458_/Y _3443_/X vssd1 vssd1 vccd1 vccd1 _3459_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_76_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6178_ _6178_/A _6178_/B vssd1 vssd1 vccd1 vccd1 _6180_/B sky130_fd_sc_hd__or2_1
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5129_ _4932_/A _4932_/B _4935_/Y _4936_/Y vssd1 vssd1 vccd1 vccd1 _5130_/C sky130_fd_sc_hd__a22oi_4
XFILLER_72_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5480_ _5634_/A vssd1 vssd1 vccd1 vccd1 _5480_/Y sky130_fd_sc_hd__inv_2
X_4500_ _4224_/C _4313_/C _4313_/B vssd1 vssd1 vccd1 vccd1 _4502_/C sky130_fd_sc_hd__a21bo_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4431_ _4569_/A vssd1 vssd1 vccd1 vccd1 _5397_/B sky130_fd_sc_hd__buf_4
XANTENNA_1 _5066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4362_ _4680_/A _4362_/B _4362_/C _5718_/A vssd1 vssd1 vccd1 vccd1 _4362_/X sky130_fd_sc_hd__and4_1
X_6101_ _6101_/A _6101_/B vssd1 vssd1 vccd1 vccd1 _6104_/C sky130_fd_sc_hd__nand2_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _4100_/A _4100_/C _4100_/B vssd1 vssd1 vccd1 vccd1 _4295_/B sky130_fd_sc_hd__a21boi_1
X_3313_ _3394_/B _3394_/C vssd1 vssd1 vccd1 vccd1 _3598_/B sky130_fd_sc_hd__nand2_2
X_6032_ _6030_/B _6030_/A _6022_/Y _6024_/Y vssd1 vssd1 vccd1 vccd1 _6037_/A sky130_fd_sc_hd__o2bb2ai_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _3246_/A _3246_/B vssd1 vssd1 vccd1 vccd1 _3245_/B sky130_fd_sc_hd__xor2_4
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ _3639_/B vssd1 vssd1 vccd1 vccd1 _3829_/B sky130_fd_sc_hd__clkbuf_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5816_ _5816_/A _5816_/B _5945_/A vssd1 vssd1 vccd1 vccd1 _5818_/B sky130_fd_sc_hd__nand3_1
X_5747_ _5742_/Y _5786_/A _5786_/B vssd1 vssd1 vccd1 vccd1 _5747_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5678_ _5678_/A _5678_/B _6127_/C _6127_/D vssd1 vssd1 vccd1 vccd1 _5840_/B sky130_fd_sc_hd__and4_2
X_4629_ _4630_/A _4630_/B _4635_/A _4635_/B vssd1 vssd1 vccd1 vccd1 _4631_/A sky130_fd_sc_hd__a22o_1
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput60 _6290_/Y vssd1 vssd1 vccd1 vccd1 r[32] sky130_fd_sc_hd__buf_2
XFILLER_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4980_ _4981_/B _4981_/C _4981_/A vssd1 vssd1 vccd1 vccd1 _4980_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3931_ _3752_/X _3757_/X _3809_/B _3809_/A vssd1 vssd1 vccd1 vccd1 _3931_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_44_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3862_ _3691_/X _3824_/Y _3829_/X _3830_/Y vssd1 vssd1 vccd1 vccd1 _3991_/A sky130_fd_sc_hd__a211o_1
X_5601_ _5592_/Y _5595_/X _5600_/Y vssd1 vssd1 vccd1 vccd1 _5601_/Y sky130_fd_sc_hd__o21ai_2
X_3793_ _3714_/X _3784_/Y _3791_/Y _3792_/X vssd1 vssd1 vccd1 vccd1 _3793_/Y sky130_fd_sc_hd__o211ai_4
X_5532_ _5532_/A _5546_/A _5532_/C _5532_/D vssd1 vssd1 vccd1 vccd1 _5532_/X sky130_fd_sc_hd__and4_1
XFILLER_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5463_ _5718_/A vssd1 vssd1 vccd1 vccd1 _5933_/D sky130_fd_sc_hd__clkbuf_2
X_5394_ _5370_/X _5371_/Y _5393_/Y vssd1 vssd1 vccd1 vccd1 _5430_/A sky130_fd_sc_hd__o21ai_4
X_4414_ _4414_/A vssd1 vssd1 vccd1 vccd1 _4414_/X sky130_fd_sc_hd__buf_2
X_4345_ _6233_/B vssd1 vssd1 vccd1 vccd1 _5348_/D sky130_fd_sc_hd__buf_2
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4276_ _4571_/A _4571_/B _5539_/B _4753_/D vssd1 vssd1 vccd1 vccd1 _4277_/B sky130_fd_sc_hd__nand4_2
X_6015_ _6023_/B vssd1 vssd1 vccd1 vccd1 _6091_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3227_ _3230_/C _3227_/B _3227_/C vssd1 vssd1 vccd1 vccd1 _3240_/A sky130_fd_sc_hd__nand3b_2
XFILLER_27_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3158_ _5229_/A vssd1 vssd1 vccd1 vccd1 _5087_/C sky130_fd_sc_hd__buf_2
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4130_ _4130_/A _4130_/B vssd1 vssd1 vccd1 vccd1 _4130_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4061_ _4906_/B vssd1 vssd1 vccd1 vccd1 _5206_/A sky130_fd_sc_hd__buf_2
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4963_ _4988_/C vssd1 vssd1 vccd1 vccd1 _5175_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3914_ _4930_/A vssd1 vssd1 vccd1 vccd1 _4619_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4894_ _4894_/A vssd1 vssd1 vccd1 vccd1 _4981_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3845_ _3845_/A _3845_/B vssd1 vssd1 vccd1 vccd1 _3999_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3776_ _3448_/A _4460_/A _3814_/A vssd1 vssd1 vccd1 vccd1 _3776_/Y sky130_fd_sc_hd__o21ai_1
X_5515_ _5515_/A _5515_/B _5515_/C vssd1 vssd1 vccd1 vccd1 _5776_/B sky130_fd_sc_hd__nand3_1
X_5446_ _5446_/A vssd1 vssd1 vccd1 vccd1 _6236_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5377_ _5372_/Y _5375_/Y _5390_/A _6202_/B vssd1 vssd1 vccd1 vccd1 _5383_/A sky130_fd_sc_hd__o2bb2ai_1
X_4328_ _4170_/X _4171_/X _4326_/Y _4327_/X vssd1 vssd1 vccd1 vccd1 _4519_/A sky130_fd_sc_hd__o211ai_2
XFILLER_59_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4259_ _4071_/A _4057_/X _4059_/Y vssd1 vssd1 vccd1 vccd1 _4259_/X sky130_fd_sc_hd__o21a_1
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3630_ _3806_/A _3630_/B _4186_/A _5834_/A vssd1 vssd1 vccd1 vccd1 _3632_/B sky130_fd_sc_hd__nand4_1
X_3561_ _3561_/A _3702_/A _3702_/B vssd1 vssd1 vccd1 vccd1 _3577_/B sky130_fd_sc_hd__nand3_2
X_5300_ _4238_/C _5299_/C _4384_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _5511_/A sky130_fd_sc_hd__a22o_2
X_6280_ _6262_/X _6258_/X _6259_/X _6258_/B _6258_/C vssd1 vssd1 vccd1 vccd1 _6285_/A
+ sky130_fd_sc_hd__a32o_1
X_3492_ _5397_/A vssd1 vssd1 vccd1 vccd1 _5580_/A sky130_fd_sc_hd__buf_4
X_5231_ _5231_/A _5378_/B vssd1 vssd1 vccd1 vccd1 _5232_/B sky130_fd_sc_hd__nand2_1
X_5162_ _4942_/Y _4943_/X _4938_/Y _4948_/Y vssd1 vssd1 vccd1 vccd1 _5163_/C sky130_fd_sc_hd__o31a_1
X_4113_ _4302_/A _4105_/B _4110_/Y vssd1 vssd1 vccd1 vccd1 _4113_/X sky130_fd_sc_hd__a21o_1
X_5093_ _5067_/A _5067_/B _5070_/A vssd1 vssd1 vccd1 vccd1 _5093_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4044_ _4044_/A vssd1 vssd1 vccd1 vccd1 _4054_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5995_ _5852_/C _6203_/D _6165_/D _5994_/A vssd1 vssd1 vccd1 vccd1 _5996_/B sky130_fd_sc_hd__a22oi_2
XFILLER_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4946_ _4933_/X _4935_/Y _4945_/X vssd1 vssd1 vccd1 vccd1 _4946_/Y sky130_fd_sc_hd__a21oi_2
X_4877_ _4877_/A _4877_/B _5207_/B _4877_/D vssd1 vssd1 vccd1 vccd1 _4878_/A sky130_fd_sc_hd__nand4_2
X_3828_ _6124_/A vssd1 vssd1 vccd1 vccd1 _6165_/A sky130_fd_sc_hd__buf_2
X_3759_ _3747_/A _3747_/B _3758_/Y vssd1 vssd1 vccd1 vccd1 _3759_/Y sky130_fd_sc_hd__o21ai_1
X_5429_ _5489_/A _5429_/B vssd1 vssd1 vccd1 vccd1 _5431_/C sky130_fd_sc_hd__nand2_1
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4800_ _4796_/A _4796_/B _4801_/A _4801_/B vssd1 vssd1 vccd1 vccd1 _4803_/B sky130_fd_sc_hd__o211ai_1
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5780_ _5780_/A _5780_/B vssd1 vssd1 vccd1 vccd1 _5780_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4731_ _4731_/A _4860_/A vssd1 vssd1 vccd1 vccd1 _4746_/A sky130_fd_sc_hd__nand2_2
X_4662_ _4399_/A _4399_/B _4394_/X _4400_/B vssd1 vssd1 vccd1 vccd1 _4669_/A sky130_fd_sc_hd__o31a_1
X_3613_ _4025_/A _5211_/A vssd1 vssd1 vccd1 vccd1 _3616_/A sky130_fd_sc_hd__nand2_1
X_4593_ _4593_/A _5223_/A vssd1 vssd1 vccd1 vccd1 _4593_/Y sky130_fd_sc_hd__nand2_1
X_3544_ _3564_/A _3564_/B _3564_/C vssd1 vssd1 vccd1 vccd1 _3565_/A sky130_fd_sc_hd__a21o_1
X_6263_ _6258_/X _6259_/X _6260_/X _6262_/X vssd1 vssd1 vccd1 vccd1 _6264_/B sky130_fd_sc_hd__a31o_1
X_3475_ _3473_/Y _5867_/A _3368_/Y _3369_/Y vssd1 vssd1 vccd1 vccd1 _3475_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5214_ _5204_/Y _5205_/X _5210_/Y _5213_/X vssd1 vssd1 vccd1 vccd1 _5222_/A sky130_fd_sc_hd__o22ai_2
X_6194_ _6119_/Y _6121_/Y _6156_/Y _6157_/X vssd1 vssd1 vccd1 vccd1 _6194_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5145_ _5145_/A vssd1 vssd1 vccd1 vccd1 _5336_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5076_ _4871_/X _5075_/Y _4865_/Y vssd1 vssd1 vccd1 vccd1 _5084_/B sky130_fd_sc_hd__a21boi_1
XFILLER_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4027_ _4025_/Y _4182_/A _4186_/A _4186_/B _4020_/Y vssd1 vssd1 vccd1 vccd1 _4177_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _5975_/B _5778_/X _5977_/Y vssd1 vssd1 vccd1 vccd1 _5978_/Y sky130_fd_sc_hd__o21bai_1
X_4929_ _4533_/X _4928_/X _4700_/Y vssd1 vssd1 vccd1 vccd1 _4929_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3322_/A vssd1 vssd1 vccd1 vccd1 _4460_/A sky130_fd_sc_hd__clkinv_4
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _3186_/X _5603_/A _3167_/Y _3190_/Y vssd1 vssd1 vccd1 vccd1 _3242_/C sky130_fd_sc_hd__o31ai_2
XFILLER_93_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5901_ _5877_/X _5869_/Y _5900_/Y vssd1 vssd1 vccd1 vccd1 _5960_/A sky130_fd_sc_hd__o21ai_1
X_5832_ _5832_/A _5832_/B vssd1 vssd1 vccd1 vccd1 _5846_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5763_ _5884_/A _5766_/B _5766_/C vssd1 vssd1 vccd1 vccd1 _5763_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_61_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4714_ _4714_/A _5134_/B vssd1 vssd1 vccd1 vccd1 _4714_/X sky130_fd_sc_hd__and2_1
X_5694_ _5694_/A _5694_/B _5694_/C vssd1 vssd1 vccd1 vccd1 _5694_/X sky130_fd_sc_hd__and3_1
X_4645_ _4645_/A _4645_/B _4645_/C vssd1 vssd1 vccd1 vccd1 _4645_/Y sky130_fd_sc_hd__nand3_2
X_4576_ _4576_/A _4576_/B _4576_/C vssd1 vssd1 vccd1 vccd1 _4605_/C sky130_fd_sc_hd__nand3_2
X_3527_ _3542_/A vssd1 vssd1 vccd1 vccd1 _4417_/A sky130_fd_sc_hd__inv_2
X_6246_ _6247_/B _6247_/A vssd1 vssd1 vccd1 vccd1 _6248_/A sky130_fd_sc_hd__nor2_1
X_3458_ _3458_/A _3458_/B _5132_/B _4625_/A vssd1 vssd1 vccd1 vccd1 _3458_/Y sky130_fd_sc_hd__nand4_4
X_6177_ _6240_/D _6240_/C _6240_/B vssd1 vssd1 vccd1 vccd1 _6178_/B sky130_fd_sc_hd__and3_1
XFILLER_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3389_ _3389_/A _3487_/A vssd1 vssd1 vccd1 vccd1 _3483_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5128_ _5128_/A _5128_/B _5299_/B _5704_/B vssd1 vssd1 vccd1 vccd1 _5130_/B sky130_fd_sc_hd__nand4_2
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5059_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5658_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_2 _5931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4430_ _4430_/A vssd1 vssd1 vccd1 vccd1 _4734_/B sky130_fd_sc_hd__buf_4
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6100_ _6151_/A _6100_/B vssd1 vssd1 vccd1 vccd1 _6101_/B sky130_fd_sc_hd__nand2_1
X_4361_ _5134_/B vssd1 vssd1 vccd1 vccd1 _5718_/A sky130_fd_sc_hd__clkbuf_4
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ _4272_/A _4294_/B _4294_/C vssd1 vssd1 vccd1 vccd1 _4295_/A sky130_fd_sc_hd__a21o_1
X_3312_ _3312_/A _3392_/A _3312_/C vssd1 vssd1 vccd1 vccd1 _3394_/C sky130_fd_sc_hd__nand3_1
X_6031_ _6022_/Y _6024_/Y _6037_/B _6030_/Y vssd1 vssd1 vccd1 vccd1 _6035_/B sky130_fd_sc_hd__o211ai_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _3199_/A _3310_/C _3310_/A _3242_/X vssd1 vssd1 vccd1 vccd1 _3246_/B sky130_fd_sc_hd__a31oi_4
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3174_ _4201_/A vssd1 vssd1 vccd1 vccd1 _3639_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5815_ _5806_/X _5807_/Y _5812_/X vssd1 vssd1 vccd1 vccd1 _5816_/A sky130_fd_sc_hd__a21o_1
X_5746_ _5732_/Y _5740_/X _5745_/X vssd1 vssd1 vccd1 vccd1 _5746_/Y sky130_fd_sc_hd__o21ai_1
X_5677_ _5677_/A vssd1 vssd1 vccd1 vccd1 _6127_/D sky130_fd_sc_hd__buf_2
X_4628_ _4628_/A _4628_/B _4628_/C vssd1 vssd1 vccd1 vccd1 _4635_/B sky130_fd_sc_hd__nand3_2
X_4559_ _4559_/A _4559_/B _4559_/C vssd1 vssd1 vccd1 vccd1 _4560_/A sky130_fd_sc_hd__nand3_1
XFILLER_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6229_ _6183_/A _6240_/A _6228_/Y _6213_/A vssd1 vssd1 vccd1 vccd1 _6230_/A sky130_fd_sc_hd__a22o_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput50 _5897_/Y vssd1 vssd1 vccd1 vccd1 r[23] sky130_fd_sc_hd__buf_2
Xoutput61 _6292_/Y vssd1 vssd1 vccd1 vccd1 r[33] sky130_fd_sc_hd__buf_2
XFILLER_68_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3930_ _3780_/X _3778_/A _3819_/B vssd1 vssd1 vccd1 vccd1 _3930_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3861_ _3859_/A _3859_/B _3860_/X _3998_/A vssd1 vssd1 vccd1 vccd1 _4005_/A sky130_fd_sc_hd__a2bb2o_1
X_3792_ _3334_/A _5656_/A _3791_/A _3790_/A vssd1 vssd1 vccd1 vccd1 _3792_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5600_ _5604_/B _5661_/A _5867_/A _6235_/B vssd1 vssd1 vccd1 vccd1 _5600_/Y sky130_fd_sc_hd__o2bb2ai_1
X_5531_ _5449_/A _5810_/B _5805_/B _5719_/C vssd1 vssd1 vccd1 vccd1 _5531_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5462_ _5432_/Y _5433_/Y _5458_/Y _5461_/Y vssd1 vssd1 vccd1 vccd1 _5479_/A sky130_fd_sc_hd__o211ai_4
X_5393_ _5612_/A _5612_/B vssd1 vssd1 vccd1 vccd1 _5393_/Y sky130_fd_sc_hd__nand2_1
X_4413_ _4630_/B _4405_/Y _4409_/X _4412_/X vssd1 vssd1 vccd1 vccd1 _4414_/A sky130_fd_sc_hd__o211ai_1
X_4344_ _6170_/B vssd1 vssd1 vccd1 vccd1 _6233_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6014_ _6011_/X _6012_/Y _6007_/X _6013_/X vssd1 vssd1 vccd1 vccd1 _6023_/B sky130_fd_sc_hd__o211ai_2
X_4275_ _4275_/A vssd1 vssd1 vccd1 vccd1 _4753_/D sky130_fd_sc_hd__buf_2
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3226_ _3226_/A _3229_/A vssd1 vssd1 vccd1 vccd1 _3227_/C sky130_fd_sc_hd__nand2_1
X_3157_ _3908_/A vssd1 vssd1 vccd1 vccd1 _5229_/A sky130_fd_sc_hd__buf_2
XFILLER_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5729_ _5729_/A _5729_/B vssd1 vssd1 vccd1 vccd1 _5730_/B sky130_fd_sc_hd__nor2_1
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4060_ _4071_/A _4057_/X _4059_/Y vssd1 vssd1 vccd1 vccd1 _4060_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4962_ _4938_/Y _4949_/Y _4951_/Y _4961_/X vssd1 vssd1 vccd1 vccd1 _4988_/C sky130_fd_sc_hd__o211ai_2
X_3913_ _3927_/A _4128_/A _4128_/B vssd1 vssd1 vccd1 vccd1 _3920_/B sky130_fd_sc_hd__nand3_1
X_4893_ _4893_/A _4893_/B _4893_/C vssd1 vssd1 vccd1 vccd1 _4894_/A sky130_fd_sc_hd__nand3_1
X_3844_ _3844_/A _3844_/B _3844_/C vssd1 vssd1 vccd1 vccd1 _3845_/A sky130_fd_sc_hd__nand3_1
X_3775_ _3679_/Y _3773_/Y _3902_/A _3676_/B vssd1 vssd1 vccd1 vccd1 _3814_/A sky130_fd_sc_hd__o2bb2ai_1
X_5514_ _5514_/A _5514_/B _5514_/C _5643_/A vssd1 vssd1 vccd1 vccd1 _5515_/C sky130_fd_sc_hd__nand4_1
X_5445_ _5445_/A _5538_/A vssd1 vssd1 vccd1 vccd1 _5445_/Y sky130_fd_sc_hd__nand2_1
X_5376_ _5376_/A vssd1 vssd1 vccd1 vccd1 _6202_/B sky130_fd_sc_hd__buf_4
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4327_ _4333_/A _4333_/B _4331_/B vssd1 vssd1 vccd1 vccd1 _4327_/X sky130_fd_sc_hd__a21o_1
X_4258_ _4088_/Y _4257_/Y _4593_/A _4619_/B _4254_/Y vssd1 vssd1 vccd1 vccd1 _4298_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3209_ _5240_/A vssd1 vssd1 vccd1 vccd1 _3458_/B sky130_fd_sc_hd__clkbuf_4
X_4189_ _3803_/B _5917_/A _5442_/C _3334_/A vssd1 vssd1 vccd1 vccd1 _4189_/Y sky130_fd_sc_hd__a22oi_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3560_ _3560_/A _3560_/B vssd1 vssd1 vccd1 vccd1 _3702_/B sky130_fd_sc_hd__nand2_1
X_3491_ _4779_/B vssd1 vssd1 vccd1 vccd1 _5578_/A sky130_fd_sc_hd__clkbuf_8
X_5230_ _5230_/A vssd1 vssd1 vccd1 vccd1 _5378_/B sky130_fd_sc_hd__buf_2
X_5161_ _5336_/A _5163_/B _5152_/X _4965_/X vssd1 vssd1 vccd1 vccd1 _5161_/X sky130_fd_sc_hd__o2bb2a_1
X_4112_ _3918_/A _3918_/C _3915_/Y vssd1 vssd1 vccd1 vccd1 _4112_/X sky130_fd_sc_hd__a21o_1
X_5092_ _5378_/A _5570_/A vssd1 vssd1 vccd1 vccd1 _5250_/A sky130_fd_sc_hd__nand2_2
X_4043_ _4043_/A _4043_/B _4043_/C vssd1 vssd1 vccd1 vccd1 _4044_/A sky130_fd_sc_hd__nand3_1
XFILLER_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5994_ _5994_/A _5994_/B _6065_/D _6165_/D vssd1 vssd1 vccd1 vccd1 _6143_/C sky130_fd_sc_hd__and4_2
X_4945_ _4945_/A _5288_/B vssd1 vssd1 vccd1 vccd1 _4945_/X sky130_fd_sc_hd__and2_1
XFILLER_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4876_ _4876_/A vssd1 vssd1 vccd1 vccd1 _4885_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3827_ _4363_/D vssd1 vssd1 vccd1 vccd1 _6124_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3758_ _3908_/A _3758_/B vssd1 vssd1 vccd1 vccd1 _3758_/Y sky130_fd_sc_hd__nand2_1
X_3689_ _3689_/A _3699_/B vssd1 vssd1 vccd1 vccd1 _3689_/Y sky130_fd_sc_hd__nand2_1
X_5428_ _5430_/A _5614_/A vssd1 vssd1 vccd1 vccd1 _5489_/A sky130_fd_sc_hd__nand2_1
X_5359_ _5513_/A _5364_/A _5364_/B vssd1 vssd1 vccd1 vccd1 _5519_/C sky130_fd_sc_hd__nand3_1
XFILLER_87_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4730_ _4730_/A _4732_/A vssd1 vssd1 vccd1 vccd1 _4860_/A sky130_fd_sc_hd__nand2_1
X_4661_ _4661_/A _4661_/B _4661_/C vssd1 vssd1 vccd1 vccd1 _4663_/B sky130_fd_sc_hd__nand3_4
XFILLER_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3612_ _3552_/A _3611_/X _3554_/Y _3555_/Y vssd1 vssd1 vccd1 vccd1 _3625_/A sky130_fd_sc_hd__a22o_1
X_4592_ _4592_/A _4592_/B vssd1 vssd1 vccd1 vccd1 _4592_/Y sky130_fd_sc_hd__nor2_1
X_3543_ _4277_/C _3543_/B vssd1 vssd1 vccd1 vccd1 _3564_/C sky130_fd_sc_hd__and2_1
X_6262_ _5506_/X _5967_/X _6255_/C _6283_/B _6235_/Y vssd1 vssd1 vccd1 vccd1 _6262_/X
+ sky130_fd_sc_hd__a41o_1
X_3474_ _3474_/A vssd1 vssd1 vccd1 vccd1 _5867_/A sky130_fd_sc_hd__clkbuf_4
X_6193_ _6193_/A _6193_/B _6193_/C vssd1 vssd1 vccd1 vccd1 _6193_/Y sky130_fd_sc_hd__nor3_1
X_5213_ _5025_/B _5403_/A _5212_/X _5208_/Y vssd1 vssd1 vccd1 vccd1 _5213_/X sky130_fd_sc_hd__o211a_2
X_5144_ _5139_/Y _5142_/X _5143_/Y vssd1 vssd1 vccd1 vccd1 _5145_/A sky130_fd_sc_hd__o21ai_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5075_ _5075_/A _5075_/B vssd1 vssd1 vccd1 vccd1 _5075_/Y sky130_fd_sc_hd__nand2_1
X_4026_ _4026_/A _5539_/A vssd1 vssd1 vccd1 vccd1 _4182_/A sky130_fd_sc_hd__nand2_4
XFILLER_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5977_ _5974_/A _5976_/Y _5974_/C vssd1 vssd1 vccd1 vccd1 _5977_/Y sky130_fd_sc_hd__o21ai_1
X_4928_ _4928_/A vssd1 vssd1 vccd1 vccd1 _4928_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_60_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4859_ _4745_/A _4858_/Y _4746_/B vssd1 vssd1 vccd1 vccd1 _5088_/B sky130_fd_sc_hd__o21ai_1
XFILLER_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _3190_/A _4827_/A _3190_/C _3829_/B vssd1 vssd1 vccd1 vccd1 _3190_/Y sky130_fd_sc_hd__nand4_1
XFILLER_66_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5900_ _5821_/A _5829_/X _5859_/Y _5863_/X vssd1 vssd1 vccd1 vccd1 _5900_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5831_ _5831_/A _5831_/B vssd1 vssd1 vccd1 vccd1 _5832_/B sky130_fd_sc_hd__nand2_1
X_5762_ _5567_/A _5567_/C _5567_/B vssd1 vssd1 vccd1 vccd1 _5766_/C sky130_fd_sc_hd__a21boi_4
XFILLER_34_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4713_ input4/X vssd1 vssd1 vccd1 vccd1 _5436_/B sky130_fd_sc_hd__clkbuf_2
X_5693_ _5672_/X _5685_/X _5744_/A _5743_/A vssd1 vssd1 vccd1 vccd1 _5693_/X sky130_fd_sc_hd__o211a_1
X_4644_ _4643_/A _4643_/B _4634_/Y _4635_/X vssd1 vssd1 vccd1 vccd1 _4645_/C sky130_fd_sc_hd__o2bb2ai_1
X_4575_ _4734_/B _4753_/D _5065_/B _5048_/A vssd1 vssd1 vccd1 vccd1 _4575_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3526_ _3342_/B _3530_/A _3461_/Y vssd1 vssd1 vccd1 vccd1 _3526_/X sky130_fd_sc_hd__o21a_1
X_6245_ _6266_/A _6245_/B vssd1 vssd1 vccd1 vccd1 _6247_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3457_ _4229_/B vssd1 vssd1 vccd1 vccd1 _4625_/A sky130_fd_sc_hd__clkbuf_4
X_6176_ _6240_/C _6240_/B _6240_/D vssd1 vssd1 vccd1 vccd1 _6178_/A sky130_fd_sc_hd__a21oi_1
X_3388_ _3388_/A _3388_/B _3388_/C vssd1 vssd1 vccd1 vccd1 _3394_/D sky130_fd_sc_hd__nand3_2
X_5127_ _4238_/C _5288_/B _5128_/A _5128_/B vssd1 vssd1 vccd1 vccd1 _5130_/A sky130_fd_sc_hd__a22o_1
X_5058_ _3189_/A _5599_/A _4853_/B _5232_/A _5081_/A vssd1 vssd1 vccd1 vccd1 _5062_/B
+ sky130_fd_sc_hd__o221ai_4
XFILLER_84_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4009_ _3938_/A _3938_/B _4133_/A _3984_/C vssd1 vssd1 vccd1 vccd1 _4009_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_44_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_3 _5534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4360_ input6/X vssd1 vssd1 vccd1 vccd1 _5134_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3311_ _3312_/A _3392_/A _3312_/C vssd1 vssd1 vccd1 vccd1 _3394_/B sky130_fd_sc_hd__a21o_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _4294_/C _4283_/Y _4284_/X _4290_/Y vssd1 vssd1 vccd1 vccd1 _4291_/Y sky130_fd_sc_hd__o2bb2ai_2
X_6030_ _6030_/A _6030_/B vssd1 vssd1 vccd1 vccd1 _6030_/Y sky130_fd_sc_hd__nand2_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _3242_/A _3242_/B _3242_/C vssd1 vssd1 vccd1 vccd1 _3242_/X sky130_fd_sc_hd__and3_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _3473_/A vssd1 vssd1 vccd1 vccd1 _4201_/A sky130_fd_sc_hd__clkbuf_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5814_ _5814_/A _5944_/A vssd1 vssd1 vccd1 vccd1 _5818_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5745_ _5742_/Y _5786_/A _5786_/B vssd1 vssd1 vccd1 vccd1 _5745_/X sky130_fd_sc_hd__a21o_1
X_5676_ _5676_/A vssd1 vssd1 vccd1 vccd1 _6127_/C sky130_fd_sc_hd__clkbuf_2
X_4627_ _3669_/X _3797_/X _4621_/A _4621_/B vssd1 vssd1 vccd1 vccd1 _4628_/C sky130_fd_sc_hd__o211ai_4
X_4558_ _4558_/A _4689_/B vssd1 vssd1 vccd1 vccd1 _4559_/C sky130_fd_sc_hd__nand2_1
X_4489_ _4489_/A _4489_/B _4489_/C _4641_/B vssd1 vssd1 vccd1 vccd1 _4490_/C sky130_fd_sc_hd__nand4_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3509_ _3509_/A _3509_/B _3509_/C vssd1 vssd1 vccd1 vccd1 _3730_/A sky130_fd_sc_hd__nand3_4
X_6228_ _6228_/A vssd1 vssd1 vccd1 vccd1 _6228_/Y sky130_fd_sc_hd__inv_2
X_6159_ _6159_/A _6159_/B vssd1 vssd1 vccd1 vccd1 _6159_/Y sky130_fd_sc_hd__nand2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput40 _4524_/X vssd1 vssd1 vccd1 vccd1 r[14] sky130_fd_sc_hd__buf_2
Xoutput51 _5982_/Y vssd1 vssd1 vccd1 vccd1 r[24] sky130_fd_sc_hd__buf_2
XFILLER_68_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput62 _3202_/Y vssd1 vssd1 vccd1 vccd1 r[3] sky130_fd_sc_hd__buf_2
XFILLER_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3860_ _3840_/X _3996_/B _3853_/Y _3849_/Y vssd1 vssd1 vccd1 vccd1 _3860_/X sky130_fd_sc_hd__o211a_1
XFILLER_31_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3791_ _3791_/A _3791_/B _3791_/C _5834_/A vssd1 vssd1 vccd1 vccd1 _3791_/Y sky130_fd_sc_hd__nand4_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5530_ _5530_/A vssd1 vssd1 vccd1 vccd1 _5719_/C sky130_fd_sc_hd__buf_2
XFILLER_31_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5461_ _5461_/A _5461_/B vssd1 vssd1 vccd1 vccd1 _5461_/Y sky130_fd_sc_hd__nand2_1
X_4412_ _4410_/Y _4630_/A _4402_/Y vssd1 vssd1 vccd1 vccd1 _4412_/X sky130_fd_sc_hd__a21o_1
X_5392_ _6236_/B _5387_/X _5388_/Y _5391_/Y vssd1 vssd1 vccd1 vccd1 _5612_/B sky130_fd_sc_hd__o211ai_4
X_4343_ _5809_/B vssd1 vssd1 vccd1 vccd1 _6170_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4274_ _4590_/B vssd1 vssd1 vccd1 vccd1 _5539_/B sky130_fd_sc_hd__clkbuf_4
X_6013_ _6165_/B _6134_/C _6006_/D _6006_/A vssd1 vssd1 vccd1 vccd1 _6013_/X sky130_fd_sc_hd__a22o_1
X_3225_ _3215_/A _3215_/B _3223_/Y vssd1 vssd1 vccd1 vccd1 _3226_/A sky130_fd_sc_hd__o21a_1
XFILLER_67_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3156_ input8/X vssd1 vssd1 vccd1 vccd1 _3908_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5728_ _5728_/A _5728_/B vssd1 vssd1 vccd1 vccd1 _5730_/A sky130_fd_sc_hd__nand2_1
X_3989_ _3837_/B _3987_/X _3988_/Y vssd1 vssd1 vccd1 vccd1 _3990_/C sky130_fd_sc_hd__o21ai_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5659_ _5833_/B _6001_/C _6003_/B _5833_/A vssd1 vssd1 vccd1 vccd1 _5659_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_89_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4961_ _4954_/Y _4948_/Y _4960_/Y vssd1 vssd1 vccd1 vccd1 _4961_/X sky130_fd_sc_hd__a21o_1
X_3912_ _3912_/A vssd1 vssd1 vccd1 vccd1 _4128_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4892_ _4768_/Y _4769_/Y _4891_/Y _4742_/A vssd1 vssd1 vccd1 vccd1 _4893_/C sky130_fd_sc_hd__a2bb2oi_2
X_3843_ _3993_/A _3833_/B _3839_/B _3839_/C vssd1 vssd1 vccd1 vccd1 _3844_/C sky130_fd_sc_hd__o211ai_1
XFILLER_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3774_ _4877_/B _3774_/B vssd1 vssd1 vccd1 vccd1 _3902_/A sky130_fd_sc_hd__nand2_2
X_5513_ _5513_/A _5513_/B vssd1 vssd1 vccd1 vccd1 _5515_/B sky130_fd_sc_hd__nand2_1
X_5444_ _5541_/A _5448_/B vssd1 vssd1 vccd1 vccd1 _5538_/A sky130_fd_sc_hd__nand2_1
X_5375_ _5375_/A _5375_/B vssd1 vssd1 vccd1 vccd1 _5375_/Y sky130_fd_sc_hd__nand2_2
XFILLER_86_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4326_ _4333_/A _4333_/B _4331_/B vssd1 vssd1 vccd1 vccd1 _4326_/Y sky130_fd_sc_hd__nand3_1
X_4257_ _4873_/A _5286_/B vssd1 vssd1 vccd1 vccd1 _4257_/Y sky130_fd_sc_hd__nand2_2
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3208_ _4738_/A vssd1 vssd1 vccd1 vccd1 _5240_/A sky130_fd_sc_hd__buf_2
X_4188_ _4530_/C vssd1 vssd1 vccd1 vccd1 _5917_/A sky130_fd_sc_hd__buf_4
XFILLER_27_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3139_ _3190_/A _4042_/B vssd1 vssd1 vccd1 vccd1 _3140_/A sky130_fd_sc_hd__and2_1
XFILLER_27_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3490_ _5212_/A vssd1 vssd1 vccd1 vccd1 _4779_/B sky130_fd_sc_hd__clkbuf_4
X_5160_ _4989_/Y _4972_/Y _4927_/Y vssd1 vssd1 vccd1 vccd1 _5178_/A sky130_fd_sc_hd__a21o_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4111_ _4103_/A _4103_/B _4110_/Y vssd1 vssd1 vccd1 vccd1 _4302_/B sky130_fd_sc_hd__o21ai_2
X_5091_ _4890_/C _5925_/B _5080_/A _5070_/C vssd1 vssd1 vccd1 vccd1 _5257_/A sky130_fd_sc_hd__a22o_1
X_4042_ _4048_/C _4042_/B _4048_/B _6203_/A vssd1 vssd1 vccd1 vccd1 _4043_/B sky130_fd_sc_hd__nand4_4
XFILLER_83_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5993_ _5948_/C _5948_/D _5992_/Y _5912_/B _5877_/X vssd1 vssd1 vccd1 vccd1 _6040_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4944_ _3448_/X _5446_/A _4533_/X _4928_/X vssd1 vssd1 vccd1 vccd1 _4944_/X sky130_fd_sc_hd__o22a_1
X_4875_ _4875_/A _4875_/B vssd1 vssd1 vccd1 vccd1 _4876_/A sky130_fd_sc_hd__nand2_1
X_3826_ _5119_/D vssd1 vssd1 vccd1 vccd1 _4363_/D sky130_fd_sc_hd__buf_4
X_3757_ _3810_/B vssd1 vssd1 vccd1 vccd1 _3757_/X sky130_fd_sc_hd__buf_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3688_ _3667_/X _3685_/B _3684_/A _3684_/B vssd1 vssd1 vccd1 vccd1 _3688_/X sky130_fd_sc_hd__o2bb2a_1
X_5427_ _5427_/A _5427_/B _5490_/A vssd1 vssd1 vccd1 vccd1 _5431_/B sky130_fd_sc_hd__nand3_1
XFILLER_87_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5358_ _5513_/A _5364_/A _5364_/B vssd1 vssd1 vccd1 vccd1 _5519_/B sky130_fd_sc_hd__a21o_1
XFILLER_59_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4309_ _4309_/A _4309_/B _4309_/C vssd1 vssd1 vccd1 vccd1 _4310_/A sky130_fd_sc_hd__nand3_1
X_5289_ _5296_/D _5296_/A _5288_/Y vssd1 vssd1 vccd1 vccd1 _5289_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_55_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _4660_/A _4660_/B vssd1 vssd1 vccd1 vccd1 _4661_/C sky130_fd_sc_hd__nand2_2
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3611_ _3611_/A vssd1 vssd1 vccd1 vccd1 _3611_/X sky130_fd_sc_hd__clkbuf_2
X_4591_ _4751_/A vssd1 vssd1 vccd1 vccd1 _4592_/B sky130_fd_sc_hd__clkbuf_2
X_3542_ _3542_/A vssd1 vssd1 vccd1 vccd1 _3543_/B sky130_fd_sc_hd__buf_2
X_6261_ _6235_/D _6235_/Y _6258_/X _6259_/X _6260_/X vssd1 vssd1 vccd1 vccd1 _6264_/A
+ sky130_fd_sc_hd__o2111ai_1
X_3473_ _3473_/A vssd1 vssd1 vccd1 vccd1 _3473_/Y sky130_fd_sc_hd__inv_2
X_6192_ _6219_/A _6219_/B _6219_/C vssd1 vssd1 vccd1 vccd1 _6193_/C sky130_fd_sc_hd__nand3_2
XFILLER_69_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5212_ _5212_/A _5212_/B vssd1 vssd1 vccd1 vccd1 _5212_/X sky130_fd_sc_hd__and2_2
XFILLER_69_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5143_ _5100_/A _5100_/B _5099_/Y vssd1 vssd1 vccd1 vccd1 _5143_/Y sky130_fd_sc_hd__a21oi_1
X_5074_ _4876_/A _4885_/C _4885_/A vssd1 vssd1 vccd1 vccd1 _5075_/B sky130_fd_sc_hd__a21o_1
XFILLER_84_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4025_ _4025_/A _5541_/A vssd1 vssd1 vccd1 vccd1 _4025_/Y sky130_fd_sc_hd__nand2_2
XFILLER_49_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5976_ _5891_/B _5891_/C _5891_/A vssd1 vssd1 vccd1 vccd1 _5976_/Y sky130_fd_sc_hd__a21oi_1
X_4927_ _4972_/A _4972_/B _4972_/C vssd1 vssd1 vccd1 vccd1 _4927_/Y sky130_fd_sc_hd__a21oi_2
X_4858_ _3533_/B _5068_/D _5245_/B _3533_/A vssd1 vssd1 vccd1 vccd1 _4858_/Y sky130_fd_sc_hd__a22oi_2
X_3809_ _3809_/A _3809_/B vssd1 vssd1 vccd1 vccd1 _3809_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4789_ _4621_/A _3795_/B _5435_/A _5449_/A _4788_/X vssd1 vssd1 vccd1 vccd1 _4950_/B
+ sky130_fd_sc_hd__a32o_2
XFILLER_87_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5830_ _3634_/X _6171_/A _5674_/B _5662_/B vssd1 vssd1 vccd1 vccd1 _5830_/X sky130_fd_sc_hd__o22a_1
XFILLER_61_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5761_ _5761_/A _5761_/B _5761_/C vssd1 vssd1 vccd1 vccd1 _5766_/B sky130_fd_sc_hd__nand3_2
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4712_ _4722_/A _4988_/A _4710_/X _4711_/Y vssd1 vssd1 vccd1 vccd1 _4712_/Y sky130_fd_sc_hd__o2bb2ai_4
X_5692_ _5840_/B _5684_/B _5672_/X _5691_/Y vssd1 vssd1 vccd1 vccd1 _5743_/A sky130_fd_sc_hd__o22ai_4
X_4643_ _4643_/A _4643_/B _4795_/A vssd1 vssd1 vccd1 vccd1 _4645_/B sky130_fd_sc_hd__nand3_1
X_4574_ _4576_/B _4576_/C _4576_/A vssd1 vssd1 vccd1 vccd1 _4574_/Y sky130_fd_sc_hd__a21oi_2
X_3525_ _3270_/B _5299_/A _4236_/B _3458_/A vssd1 vssd1 vccd1 vccd1 _3525_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6244_ _6244_/A _6244_/B _6244_/C vssd1 vssd1 vccd1 vccd1 _6245_/B sky130_fd_sc_hd__nand3_1
X_3456_ _3766_/A vssd1 vssd1 vccd1 vccd1 _4229_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_39_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6175_ _6139_/B _6139_/C _6131_/X vssd1 vssd1 vccd1 vccd1 _6240_/D sky130_fd_sc_hd__a21o_1
X_3387_ _3392_/A _3392_/D vssd1 vssd1 vccd1 vccd1 _3388_/C sky130_fd_sc_hd__nand2_1
X_5126_ _5120_/Y _5121_/Y _5122_/X _5125_/X vssd1 vssd1 vccd1 vccd1 _5126_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_57_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5057_ _4860_/X _5046_/A _4868_/Y _5051_/Y vssd1 vssd1 vccd1 vccd1 _5062_/A sky130_fd_sc_hd__o22a_1
X_4008_ _4008_/A _4008_/B _4008_/C vssd1 vssd1 vccd1 vccd1 _4008_/X sky130_fd_sc_hd__and3_1
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5959_ _5966_/C _5959_/B _5959_/C vssd1 vssd1 vccd1 vccd1 _6058_/A sky130_fd_sc_hd__nand3b_1
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_4 _4674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3310_ _3310_/A _3310_/B _3310_/C _5845_/A vssd1 vssd1 vccd1 vccd1 _3312_/C sky130_fd_sc_hd__and4_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ _4091_/A _4091_/B _4288_/Y _4289_/X vssd1 vssd1 vccd1 vccd1 _4290_/Y sky130_fd_sc_hd__a22oi_4
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3241_/A _3241_/B vssd1 vssd1 vccd1 vccd1 _3246_/A sky130_fd_sc_hd__nand2_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3172_ _3170_/A _3170_/B _6297_/A vssd1 vssd1 vccd1 vccd1 _3202_/A sky130_fd_sc_hd__o21ai_2
XFILLER_94_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5813_ _5806_/X _5807_/Y _5812_/X vssd1 vssd1 vccd1 vccd1 _5944_/A sky130_fd_sc_hd__a21oi_2
XFILLER_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5744_ _5744_/A vssd1 vssd1 vccd1 vccd1 _5786_/B sky130_fd_sc_hd__clkbuf_2
X_5675_ _5399_/Y _5580_/Y _5674_/X _5585_/A vssd1 vssd1 vccd1 vccd1 _5675_/X sky130_fd_sc_hd__a22o_2
X_4626_ _4621_/A _4621_/B _4625_/Y vssd1 vssd1 vccd1 vccd1 _4628_/B sky130_fd_sc_hd__a21o_1
X_4557_ _4557_/A _4557_/B vssd1 vssd1 vccd1 vccd1 _4558_/A sky130_fd_sc_hd__nand2_1
X_4488_ _4281_/X _4291_/Y _4308_/A _4487_/Y vssd1 vssd1 vccd1 vccd1 _4490_/B sky130_fd_sc_hd__a2bb2oi_1
X_3508_ _3641_/A _4422_/B _3514_/A _3508_/D vssd1 vssd1 vccd1 vccd1 _3509_/C sky130_fd_sc_hd__nand4_1
XFILLER_89_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6227_ _6227_/A vssd1 vssd1 vccd1 vccd1 _6240_/A sky130_fd_sc_hd__inv_2
X_3439_ _3439_/A _5132_/A _5087_/C vssd1 vssd1 vccd1 vccd1 _3445_/A sky130_fd_sc_hd__nand3_1
X_6158_ _6119_/Y _6121_/Y _6156_/Y _6157_/X vssd1 vssd1 vccd1 vccd1 _6161_/A sky130_fd_sc_hd__o211a_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5109_ _5310_/A _5309_/A _5309_/B vssd1 vssd1 vccd1 vccd1 _5110_/B sky130_fd_sc_hd__nand3_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6089_ _6089_/A _6089_/B _6089_/C vssd1 vssd1 vccd1 vccd1 _6090_/B sky130_fd_sc_hd__nand3_1
XFILLER_13_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput52 _6060_/Y vssd1 vssd1 vccd1 vccd1 r[25] sky130_fd_sc_hd__buf_2
Xoutput41 _4686_/Y vssd1 vssd1 vccd1 vccd1 r[15] sky130_fd_sc_hd__buf_2
Xoutput63 _3245_/Y vssd1 vssd1 vccd1 vccd1 r[4] sky130_fd_sc_hd__buf_2
XFILLER_95_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3790_ _3790_/A vssd1 vssd1 vccd1 vccd1 _3791_/B sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5460_ _5460_/A _5460_/B vssd1 vssd1 vccd1 vccd1 _5461_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4411_ _4411_/A _4411_/B vssd1 vssd1 vccd1 vccd1 _4630_/A sky130_fd_sc_hd__nand2_2
X_5391_ _5391_/A _5391_/B vssd1 vssd1 vccd1 vccd1 _5391_/Y sky130_fd_sc_hd__nand2_1
X_4342_ _4338_/A _4169_/X _4340_/A _4340_/B _4341_/X vssd1 vssd1 vccd1 vccd1 _4342_/X
+ sky130_fd_sc_hd__a41o_4
X_4273_ _3189_/A _4261_/Y _4270_/A vssd1 vssd1 vccd1 vccd1 _4279_/A sky130_fd_sc_hd__o21ai_1
X_3224_ _3229_/A _3229_/B _3223_/Y vssd1 vssd1 vccd1 vccd1 _3227_/B sky130_fd_sc_hd__a21o_1
X_6012_ _6127_/B _6170_/C _6170_/D _3829_/C vssd1 vssd1 vccd1 vccd1 _6012_/Y sky130_fd_sc_hd__a22oi_2
.ends

