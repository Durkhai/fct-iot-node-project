magic
tech sky130A
magscale 1 2
timestamp 1653581497
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 1980 178848 117552
<< metal2 >>
rect 1490 119200 1546 120000
rect 4434 119200 4490 120000
rect 7378 119200 7434 120000
rect 10322 119200 10378 120000
rect 13266 119200 13322 120000
rect 16210 119200 16266 120000
rect 19154 119200 19210 120000
rect 22098 119200 22154 120000
rect 25042 119200 25098 120000
rect 27986 119200 28042 120000
rect 30930 119200 30986 120000
rect 33874 119200 33930 120000
rect 36818 119200 36874 120000
rect 39854 119200 39910 120000
rect 42798 119200 42854 120000
rect 45742 119200 45798 120000
rect 48686 119200 48742 120000
rect 51630 119200 51686 120000
rect 54574 119200 54630 120000
rect 57518 119200 57574 120000
rect 60462 119200 60518 120000
rect 63406 119200 63462 120000
rect 66350 119200 66406 120000
rect 69294 119200 69350 120000
rect 72238 119200 72294 120000
rect 75274 119200 75330 120000
rect 78218 119200 78274 120000
rect 81162 119200 81218 120000
rect 84106 119200 84162 120000
rect 87050 119200 87106 120000
rect 89994 119200 90050 120000
rect 92938 119200 92994 120000
rect 95882 119200 95938 120000
rect 98826 119200 98882 120000
rect 101770 119200 101826 120000
rect 104714 119200 104770 120000
rect 107658 119200 107714 120000
rect 110694 119200 110750 120000
rect 113638 119200 113694 120000
rect 116582 119200 116638 120000
rect 119526 119200 119582 120000
rect 122470 119200 122526 120000
rect 125414 119200 125470 120000
rect 128358 119200 128414 120000
rect 131302 119200 131358 120000
rect 134246 119200 134302 120000
rect 137190 119200 137246 120000
rect 140134 119200 140190 120000
rect 143078 119200 143134 120000
rect 146114 119200 146170 120000
rect 149058 119200 149114 120000
rect 152002 119200 152058 120000
rect 154946 119200 155002 120000
rect 157890 119200 157946 120000
rect 160834 119200 160890 120000
rect 163778 119200 163834 120000
rect 166722 119200 166778 120000
rect 169666 119200 169722 120000
rect 172610 119200 172666 120000
rect 175554 119200 175610 120000
rect 178498 119200 178554 120000
rect 1398 0 1454 800
rect 4158 0 4214 800
rect 6918 0 6974 800
rect 9678 0 9734 800
rect 12438 0 12494 800
rect 15198 0 15254 800
rect 17958 0 18014 800
rect 20718 0 20774 800
rect 23478 0 23534 800
rect 26238 0 26294 800
rect 29090 0 29146 800
rect 31850 0 31906 800
rect 34610 0 34666 800
rect 37370 0 37426 800
rect 40130 0 40186 800
rect 42890 0 42946 800
rect 45650 0 45706 800
rect 48410 0 48466 800
rect 51170 0 51226 800
rect 54022 0 54078 800
rect 56782 0 56838 800
rect 59542 0 59598 800
rect 62302 0 62358 800
rect 65062 0 65118 800
rect 67822 0 67878 800
rect 70582 0 70638 800
rect 73342 0 73398 800
rect 76102 0 76158 800
rect 78954 0 79010 800
rect 81714 0 81770 800
rect 84474 0 84530 800
rect 87234 0 87290 800
rect 89994 0 90050 800
rect 92754 0 92810 800
rect 95514 0 95570 800
rect 98274 0 98330 800
rect 101034 0 101090 800
rect 103794 0 103850 800
rect 106646 0 106702 800
rect 109406 0 109462 800
rect 112166 0 112222 800
rect 114926 0 114982 800
rect 117686 0 117742 800
rect 120446 0 120502 800
rect 123206 0 123262 800
rect 125966 0 126022 800
rect 128726 0 128782 800
rect 131578 0 131634 800
rect 134338 0 134394 800
rect 137098 0 137154 800
rect 139858 0 139914 800
rect 142618 0 142674 800
rect 145378 0 145434 800
rect 148138 0 148194 800
rect 150898 0 150954 800
rect 153658 0 153714 800
rect 156510 0 156566 800
rect 159270 0 159326 800
rect 162030 0 162086 800
rect 164790 0 164846 800
rect 167550 0 167606 800
rect 170310 0 170366 800
rect 173070 0 173126 800
rect 175830 0 175886 800
rect 178590 0 178646 800
<< obsm2 >>
rect 1398 119144 1434 119354
rect 1602 119144 4378 119354
rect 4546 119144 7322 119354
rect 7490 119144 10266 119354
rect 10434 119144 13210 119354
rect 13378 119144 16154 119354
rect 16322 119144 19098 119354
rect 19266 119144 22042 119354
rect 22210 119144 24986 119354
rect 25154 119144 27930 119354
rect 28098 119144 30874 119354
rect 31042 119144 33818 119354
rect 33986 119144 36762 119354
rect 36930 119144 39798 119354
rect 39966 119144 42742 119354
rect 42910 119144 45686 119354
rect 45854 119144 48630 119354
rect 48798 119144 51574 119354
rect 51742 119144 54518 119354
rect 54686 119144 57462 119354
rect 57630 119144 60406 119354
rect 60574 119144 63350 119354
rect 63518 119144 66294 119354
rect 66462 119144 69238 119354
rect 69406 119144 72182 119354
rect 72350 119144 75218 119354
rect 75386 119144 78162 119354
rect 78330 119144 81106 119354
rect 81274 119144 84050 119354
rect 84218 119144 86994 119354
rect 87162 119144 89938 119354
rect 90106 119144 92882 119354
rect 93050 119144 95826 119354
rect 95994 119144 98770 119354
rect 98938 119144 101714 119354
rect 101882 119144 104658 119354
rect 104826 119144 107602 119354
rect 107770 119144 110638 119354
rect 110806 119144 113582 119354
rect 113750 119144 116526 119354
rect 116694 119144 119470 119354
rect 119638 119144 122414 119354
rect 122582 119144 125358 119354
rect 125526 119144 128302 119354
rect 128470 119144 131246 119354
rect 131414 119144 134190 119354
rect 134358 119144 137134 119354
rect 137302 119144 140078 119354
rect 140246 119144 143022 119354
rect 143190 119144 146058 119354
rect 146226 119144 149002 119354
rect 149170 119144 151946 119354
rect 152114 119144 154890 119354
rect 155058 119144 157834 119354
rect 158002 119144 160778 119354
rect 160946 119144 163722 119354
rect 163890 119144 166666 119354
rect 166834 119144 169610 119354
rect 169778 119144 172554 119354
rect 172722 119144 175498 119354
rect 175666 119144 178442 119354
rect 178610 119144 178644 119354
rect 1398 856 178644 119144
rect 1510 711 4102 856
rect 4270 711 6862 856
rect 7030 711 9622 856
rect 9790 711 12382 856
rect 12550 711 15142 856
rect 15310 711 17902 856
rect 18070 711 20662 856
rect 20830 711 23422 856
rect 23590 711 26182 856
rect 26350 711 29034 856
rect 29202 711 31794 856
rect 31962 711 34554 856
rect 34722 711 37314 856
rect 37482 711 40074 856
rect 40242 711 42834 856
rect 43002 711 45594 856
rect 45762 711 48354 856
rect 48522 711 51114 856
rect 51282 711 53966 856
rect 54134 711 56726 856
rect 56894 711 59486 856
rect 59654 711 62246 856
rect 62414 711 65006 856
rect 65174 711 67766 856
rect 67934 711 70526 856
rect 70694 711 73286 856
rect 73454 711 76046 856
rect 76214 711 78898 856
rect 79066 711 81658 856
rect 81826 711 84418 856
rect 84586 711 87178 856
rect 87346 711 89938 856
rect 90106 711 92698 856
rect 92866 711 95458 856
rect 95626 711 98218 856
rect 98386 711 100978 856
rect 101146 711 103738 856
rect 103906 711 106590 856
rect 106758 711 109350 856
rect 109518 711 112110 856
rect 112278 711 114870 856
rect 115038 711 117630 856
rect 117798 711 120390 856
rect 120558 711 123150 856
rect 123318 711 125910 856
rect 126078 711 128670 856
rect 128838 711 131522 856
rect 131690 711 134282 856
rect 134450 711 137042 856
rect 137210 711 139802 856
rect 139970 711 142562 856
rect 142730 711 145322 856
rect 145490 711 148082 856
rect 148250 711 150842 856
rect 151010 711 153602 856
rect 153770 711 156454 856
rect 156622 711 159214 856
rect 159382 711 161974 856
rect 162142 711 164734 856
rect 164902 711 167494 856
rect 167662 711 170254 856
rect 170422 711 173014 856
rect 173182 711 175774 856
rect 175942 711 178534 856
<< metal3 >>
rect 0 119008 800 119128
rect 179200 118872 180000 118992
rect 0 117376 800 117496
rect 179200 116968 180000 117088
rect 0 115880 800 116000
rect 179200 115064 180000 115184
rect 0 114248 800 114368
rect 179200 113160 180000 113280
rect 0 112616 800 112736
rect 179200 111392 180000 111512
rect 0 111120 800 111240
rect 0 109488 800 109608
rect 179200 109488 180000 109608
rect 0 107992 800 108112
rect 179200 107584 180000 107704
rect 0 106360 800 106480
rect 179200 105680 180000 105800
rect 0 104728 800 104848
rect 179200 103776 180000 103896
rect 0 103232 800 103352
rect 179200 102008 180000 102128
rect 0 101600 800 101720
rect 0 100104 800 100224
rect 179200 100104 180000 100224
rect 0 98472 800 98592
rect 179200 98200 180000 98320
rect 0 96840 800 96960
rect 179200 96296 180000 96416
rect 0 95344 800 95464
rect 179200 94528 180000 94648
rect 0 93712 800 93832
rect 179200 92624 180000 92744
rect 0 92216 800 92336
rect 0 90584 800 90704
rect 179200 90720 180000 90840
rect 0 88952 800 89072
rect 179200 88816 180000 88936
rect 0 87456 800 87576
rect 179200 86912 180000 87032
rect 0 85824 800 85944
rect 179200 85144 180000 85264
rect 0 84328 800 84448
rect 179200 83240 180000 83360
rect 0 82696 800 82816
rect 179200 81336 180000 81456
rect 0 81064 800 81184
rect 0 79568 800 79688
rect 179200 79432 180000 79552
rect 0 77936 800 78056
rect 179200 77664 180000 77784
rect 0 76440 800 76560
rect 179200 75760 180000 75880
rect 0 74808 800 74928
rect 179200 73856 180000 73976
rect 0 73176 800 73296
rect 179200 71952 180000 72072
rect 0 71680 800 71800
rect 0 70048 800 70168
rect 179200 70048 180000 70168
rect 0 68552 800 68672
rect 179200 68280 180000 68400
rect 0 66920 800 67040
rect 179200 66376 180000 66496
rect 0 65288 800 65408
rect 179200 64472 180000 64592
rect 0 63792 800 63912
rect 179200 62568 180000 62688
rect 0 62160 800 62280
rect 0 60664 800 60784
rect 179200 60800 180000 60920
rect 0 59032 800 59152
rect 179200 58896 180000 59016
rect 0 57400 800 57520
rect 179200 56992 180000 57112
rect 0 55904 800 56024
rect 179200 55088 180000 55208
rect 0 54272 800 54392
rect 179200 53184 180000 53304
rect 0 52640 800 52760
rect 179200 51416 180000 51536
rect 0 51144 800 51264
rect 0 49512 800 49632
rect 179200 49512 180000 49632
rect 0 48016 800 48136
rect 179200 47608 180000 47728
rect 0 46384 800 46504
rect 179200 45704 180000 45824
rect 0 44752 800 44872
rect 179200 43800 180000 43920
rect 0 43256 800 43376
rect 179200 42032 180000 42152
rect 0 41624 800 41744
rect 0 40128 800 40248
rect 179200 40128 180000 40248
rect 0 38496 800 38616
rect 179200 38224 180000 38344
rect 0 36864 800 36984
rect 179200 36320 180000 36440
rect 0 35368 800 35488
rect 179200 34552 180000 34672
rect 0 33736 800 33856
rect 179200 32648 180000 32768
rect 0 32240 800 32360
rect 0 30608 800 30728
rect 179200 30744 180000 30864
rect 0 28976 800 29096
rect 179200 28840 180000 28960
rect 0 27480 800 27600
rect 179200 26936 180000 27056
rect 0 25848 800 25968
rect 179200 25168 180000 25288
rect 0 24352 800 24472
rect 179200 23264 180000 23384
rect 0 22720 800 22840
rect 179200 21360 180000 21480
rect 0 21088 800 21208
rect 0 19592 800 19712
rect 179200 19456 180000 19576
rect 0 17960 800 18080
rect 179200 17688 180000 17808
rect 0 16464 800 16584
rect 179200 15784 180000 15904
rect 0 14832 800 14952
rect 179200 13880 180000 14000
rect 0 13200 800 13320
rect 179200 11976 180000 12096
rect 0 11704 800 11824
rect 0 10072 800 10192
rect 179200 10072 180000 10192
rect 0 8576 800 8696
rect 179200 8304 180000 8424
rect 0 6944 800 7064
rect 179200 6400 180000 6520
rect 0 5312 800 5432
rect 179200 4496 180000 4616
rect 0 3816 800 3936
rect 179200 2592 180000 2712
rect 0 2184 800 2304
rect 0 688 800 808
rect 179200 824 180000 944
<< obsm3 >>
rect 880 119072 179200 119101
rect 880 118928 179120 119072
rect 800 118792 179120 118928
rect 800 117576 179200 118792
rect 880 117296 179200 117576
rect 800 117168 179200 117296
rect 800 116888 179120 117168
rect 800 116080 179200 116888
rect 880 115800 179200 116080
rect 800 115264 179200 115800
rect 800 114984 179120 115264
rect 800 114448 179200 114984
rect 880 114168 179200 114448
rect 800 113360 179200 114168
rect 800 113080 179120 113360
rect 800 112816 179200 113080
rect 880 112536 179200 112816
rect 800 111592 179200 112536
rect 800 111320 179120 111592
rect 880 111312 179120 111320
rect 880 111040 179200 111312
rect 800 109688 179200 111040
rect 880 109408 179120 109688
rect 800 108192 179200 109408
rect 880 107912 179200 108192
rect 800 107784 179200 107912
rect 800 107504 179120 107784
rect 800 106560 179200 107504
rect 880 106280 179200 106560
rect 800 105880 179200 106280
rect 800 105600 179120 105880
rect 800 104928 179200 105600
rect 880 104648 179200 104928
rect 800 103976 179200 104648
rect 800 103696 179120 103976
rect 800 103432 179200 103696
rect 880 103152 179200 103432
rect 800 102208 179200 103152
rect 800 101928 179120 102208
rect 800 101800 179200 101928
rect 880 101520 179200 101800
rect 800 100304 179200 101520
rect 880 100024 179120 100304
rect 800 98672 179200 100024
rect 880 98400 179200 98672
rect 880 98392 179120 98400
rect 800 98120 179120 98392
rect 800 97040 179200 98120
rect 880 96760 179200 97040
rect 800 96496 179200 96760
rect 800 96216 179120 96496
rect 800 95544 179200 96216
rect 880 95264 179200 95544
rect 800 94728 179200 95264
rect 800 94448 179120 94728
rect 800 93912 179200 94448
rect 880 93632 179200 93912
rect 800 92824 179200 93632
rect 800 92544 179120 92824
rect 800 92416 179200 92544
rect 880 92136 179200 92416
rect 800 90920 179200 92136
rect 800 90784 179120 90920
rect 880 90640 179120 90784
rect 880 90504 179200 90640
rect 800 89152 179200 90504
rect 880 89016 179200 89152
rect 880 88872 179120 89016
rect 800 88736 179120 88872
rect 800 87656 179200 88736
rect 880 87376 179200 87656
rect 800 87112 179200 87376
rect 800 86832 179120 87112
rect 800 86024 179200 86832
rect 880 85744 179200 86024
rect 800 85344 179200 85744
rect 800 85064 179120 85344
rect 800 84528 179200 85064
rect 880 84248 179200 84528
rect 800 83440 179200 84248
rect 800 83160 179120 83440
rect 800 82896 179200 83160
rect 880 82616 179200 82896
rect 800 81536 179200 82616
rect 800 81264 179120 81536
rect 880 81256 179120 81264
rect 880 80984 179200 81256
rect 800 79768 179200 80984
rect 880 79632 179200 79768
rect 880 79488 179120 79632
rect 800 79352 179120 79488
rect 800 78136 179200 79352
rect 880 77864 179200 78136
rect 880 77856 179120 77864
rect 800 77584 179120 77856
rect 800 76640 179200 77584
rect 880 76360 179200 76640
rect 800 75960 179200 76360
rect 800 75680 179120 75960
rect 800 75008 179200 75680
rect 880 74728 179200 75008
rect 800 74056 179200 74728
rect 800 73776 179120 74056
rect 800 73376 179200 73776
rect 880 73096 179200 73376
rect 800 72152 179200 73096
rect 800 71880 179120 72152
rect 880 71872 179120 71880
rect 880 71600 179200 71872
rect 800 70248 179200 71600
rect 880 69968 179120 70248
rect 800 68752 179200 69968
rect 880 68480 179200 68752
rect 880 68472 179120 68480
rect 800 68200 179120 68472
rect 800 67120 179200 68200
rect 880 66840 179200 67120
rect 800 66576 179200 66840
rect 800 66296 179120 66576
rect 800 65488 179200 66296
rect 880 65208 179200 65488
rect 800 64672 179200 65208
rect 800 64392 179120 64672
rect 800 63992 179200 64392
rect 880 63712 179200 63992
rect 800 62768 179200 63712
rect 800 62488 179120 62768
rect 800 62360 179200 62488
rect 880 62080 179200 62360
rect 800 61000 179200 62080
rect 800 60864 179120 61000
rect 880 60720 179120 60864
rect 880 60584 179200 60720
rect 800 59232 179200 60584
rect 880 59096 179200 59232
rect 880 58952 179120 59096
rect 800 58816 179120 58952
rect 800 57600 179200 58816
rect 880 57320 179200 57600
rect 800 57192 179200 57320
rect 800 56912 179120 57192
rect 800 56104 179200 56912
rect 880 55824 179200 56104
rect 800 55288 179200 55824
rect 800 55008 179120 55288
rect 800 54472 179200 55008
rect 880 54192 179200 54472
rect 800 53384 179200 54192
rect 800 53104 179120 53384
rect 800 52840 179200 53104
rect 880 52560 179200 52840
rect 800 51616 179200 52560
rect 800 51344 179120 51616
rect 880 51336 179120 51344
rect 880 51064 179200 51336
rect 800 49712 179200 51064
rect 880 49432 179120 49712
rect 800 48216 179200 49432
rect 880 47936 179200 48216
rect 800 47808 179200 47936
rect 800 47528 179120 47808
rect 800 46584 179200 47528
rect 880 46304 179200 46584
rect 800 45904 179200 46304
rect 800 45624 179120 45904
rect 800 44952 179200 45624
rect 880 44672 179200 44952
rect 800 44000 179200 44672
rect 800 43720 179120 44000
rect 800 43456 179200 43720
rect 880 43176 179200 43456
rect 800 42232 179200 43176
rect 800 41952 179120 42232
rect 800 41824 179200 41952
rect 880 41544 179200 41824
rect 800 40328 179200 41544
rect 880 40048 179120 40328
rect 800 38696 179200 40048
rect 880 38424 179200 38696
rect 880 38416 179120 38424
rect 800 38144 179120 38416
rect 800 37064 179200 38144
rect 880 36784 179200 37064
rect 800 36520 179200 36784
rect 800 36240 179120 36520
rect 800 35568 179200 36240
rect 880 35288 179200 35568
rect 800 34752 179200 35288
rect 800 34472 179120 34752
rect 800 33936 179200 34472
rect 880 33656 179200 33936
rect 800 32848 179200 33656
rect 800 32568 179120 32848
rect 800 32440 179200 32568
rect 880 32160 179200 32440
rect 800 30944 179200 32160
rect 800 30808 179120 30944
rect 880 30664 179120 30808
rect 880 30528 179200 30664
rect 800 29176 179200 30528
rect 880 29040 179200 29176
rect 880 28896 179120 29040
rect 800 28760 179120 28896
rect 800 27680 179200 28760
rect 880 27400 179200 27680
rect 800 27136 179200 27400
rect 800 26856 179120 27136
rect 800 26048 179200 26856
rect 880 25768 179200 26048
rect 800 25368 179200 25768
rect 800 25088 179120 25368
rect 800 24552 179200 25088
rect 880 24272 179200 24552
rect 800 23464 179200 24272
rect 800 23184 179120 23464
rect 800 22920 179200 23184
rect 880 22640 179200 22920
rect 800 21560 179200 22640
rect 800 21288 179120 21560
rect 880 21280 179120 21288
rect 880 21008 179200 21280
rect 800 19792 179200 21008
rect 880 19656 179200 19792
rect 880 19512 179120 19656
rect 800 19376 179120 19512
rect 800 18160 179200 19376
rect 880 17888 179200 18160
rect 880 17880 179120 17888
rect 800 17608 179120 17880
rect 800 16664 179200 17608
rect 880 16384 179200 16664
rect 800 15984 179200 16384
rect 800 15704 179120 15984
rect 800 15032 179200 15704
rect 880 14752 179200 15032
rect 800 14080 179200 14752
rect 800 13800 179120 14080
rect 800 13400 179200 13800
rect 880 13120 179200 13400
rect 800 12176 179200 13120
rect 800 11904 179120 12176
rect 880 11896 179120 11904
rect 880 11624 179200 11896
rect 800 10272 179200 11624
rect 880 9992 179120 10272
rect 800 8776 179200 9992
rect 880 8504 179200 8776
rect 880 8496 179120 8504
rect 800 8224 179120 8496
rect 800 7144 179200 8224
rect 880 6864 179200 7144
rect 800 6600 179200 6864
rect 800 6320 179120 6600
rect 800 5512 179200 6320
rect 880 5232 179200 5512
rect 800 4696 179200 5232
rect 800 4416 179120 4696
rect 800 4016 179200 4416
rect 880 3736 179200 4016
rect 800 2792 179200 3736
rect 800 2512 179120 2792
rect 800 2384 179200 2512
rect 880 2104 179200 2384
rect 800 1024 179200 2104
rect 800 888 179120 1024
rect 880 744 179120 888
rect 880 715 179200 744
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 57099 3435 65568 113933
rect 66048 3435 80928 113933
rect 81408 3435 96288 113933
rect 96768 3435 111648 113933
rect 112128 3435 114757 113933
<< labels >>
rlabel metal2 s 4434 119200 4490 120000 6 a11[0]
port 1 nsew signal output
rlabel metal3 s 179200 42032 180000 42152 6 a11[10]
port 2 nsew signal output
rlabel metal2 s 63406 119200 63462 120000 6 a11[11]
port 3 nsew signal output
rlabel metal3 s 0 66920 800 67040 6 a11[12]
port 4 nsew signal output
rlabel metal3 s 179200 51416 180000 51536 6 a11[13]
port 5 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 a11[14]
port 6 nsew signal output
rlabel metal3 s 179200 60800 180000 60920 6 a11[15]
port 7 nsew signal output
rlabel metal3 s 179200 62568 180000 62688 6 a11[16]
port 8 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 a11[17]
port 9 nsew signal output
rlabel metal3 s 179200 73856 180000 73976 6 a11[18]
port 10 nsew signal output
rlabel metal3 s 0 88952 800 89072 6 a11[19]
port 11 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 a11[1]
port 12 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 a11[20]
port 13 nsew signal output
rlabel metal2 s 104714 119200 104770 120000 6 a11[21]
port 14 nsew signal output
rlabel metal3 s 0 96840 800 96960 6 a11[22]
port 15 nsew signal output
rlabel metal3 s 179200 96296 180000 96416 6 a11[23]
port 16 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 a11[24]
port 17 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 a11[25]
port 18 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 a11[26]
port 19 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 a11[27]
port 20 nsew signal output
rlabel metal3 s 179200 113160 180000 113280 6 a11[28]
port 21 nsew signal output
rlabel metal2 s 154946 119200 155002 120000 6 a11[29]
port 22 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 a11[2]
port 23 nsew signal output
rlabel metal2 s 167550 0 167606 800 6 a11[30]
port 24 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 a11[31]
port 25 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 a11[3]
port 26 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 a11[4]
port 27 nsew signal output
rlabel metal3 s 179200 26936 180000 27056 6 a11[5]
port 28 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 a11[6]
port 29 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 a11[7]
port 30 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 a11[8]
port 31 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 a11[9]
port 32 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 a12[0]
port 33 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 a12[10]
port 34 nsew signal output
rlabel metal2 s 66350 119200 66406 120000 6 a12[11]
port 35 nsew signal output
rlabel metal3 s 179200 47608 180000 47728 6 a12[12]
port 36 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 a12[13]
port 37 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 a12[14]
port 38 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 a12[15]
port 39 nsew signal output
rlabel metal3 s 179200 64472 180000 64592 6 a12[16]
port 40 nsew signal output
rlabel metal3 s 179200 68280 180000 68400 6 a12[17]
port 41 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 a12[18]
port 42 nsew signal output
rlabel metal2 s 101770 119200 101826 120000 6 a12[19]
port 43 nsew signal output
rlabel metal3 s 179200 4496 180000 4616 6 a12[1]
port 44 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 a12[20]
port 45 nsew signal output
rlabel metal3 s 179200 83240 180000 83360 6 a12[21]
port 46 nsew signal output
rlabel metal3 s 0 98472 800 98592 6 a12[22]
port 47 nsew signal output
rlabel metal3 s 0 101600 800 101720 6 a12[23]
port 48 nsew signal output
rlabel metal3 s 179200 98200 180000 98320 6 a12[24]
port 49 nsew signal output
rlabel metal3 s 179200 103776 180000 103896 6 a12[25]
port 50 nsew signal output
rlabel metal3 s 179200 107584 180000 107704 6 a12[26]
port 51 nsew signal output
rlabel metal2 s 159270 0 159326 800 6 a12[27]
port 52 nsew signal output
rlabel metal2 s 140134 119200 140190 120000 6 a12[28]
port 53 nsew signal output
rlabel metal3 s 0 112616 800 112736 6 a12[29]
port 54 nsew signal output
rlabel metal3 s 179200 10072 180000 10192 6 a12[2]
port 55 nsew signal output
rlabel metal3 s 0 114248 800 114368 6 a12[30]
port 56 nsew signal output
rlabel metal2 s 172610 119200 172666 120000 6 a12[31]
port 57 nsew signal output
rlabel metal3 s 179200 15784 180000 15904 6 a12[3]
port 58 nsew signal output
rlabel metal2 s 33874 119200 33930 120000 6 a12[4]
port 59 nsew signal output
rlabel metal3 s 0 32240 800 32360 6 a12[5]
port 60 nsew signal output
rlabel metal3 s 179200 28840 180000 28960 6 a12[6]
port 61 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 a12[7]
port 62 nsew signal output
rlabel metal3 s 0 46384 800 46504 6 a12[8]
port 63 nsew signal output
rlabel metal3 s 179200 36320 180000 36440 6 a12[9]
port 64 nsew signal output
rlabel metal2 s 1490 119200 1546 120000 6 ack_o
port 65 nsew signal output
rlabel metal2 s 7378 119200 7434 120000 6 adr_i[0]
port 66 nsew signal input
rlabel metal3 s 179200 6400 180000 6520 6 adr_i[1]
port 67 nsew signal input
rlabel metal3 s 179200 11976 180000 12096 6 adr_i[2]
port 68 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 adr_i[3]
port 69 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 b10[0]
port 70 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 b10[10]
port 71 nsew signal output
rlabel metal2 s 69294 119200 69350 120000 6 b10[11]
port 72 nsew signal output
rlabel metal3 s 0 68552 800 68672 6 b10[12]
port 73 nsew signal output
rlabel metal2 s 75274 119200 75330 120000 6 b10[13]
port 74 nsew signal output
rlabel metal2 s 78218 119200 78274 120000 6 b10[14]
port 75 nsew signal output
rlabel metal3 s 0 81064 800 81184 6 b10[15]
port 76 nsew signal output
rlabel metal2 s 87050 119200 87106 120000 6 b10[16]
port 77 nsew signal output
rlabel metal2 s 95882 119200 95938 120000 6 b10[17]
port 78 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 b10[18]
port 79 nsew signal output
rlabel metal2 s 123206 0 123262 800 6 b10[19]
port 80 nsew signal output
rlabel metal3 s 179200 8304 180000 8424 6 b10[1]
port 81 nsew signal output
rlabel metal2 s 131578 0 131634 800 6 b10[20]
port 82 nsew signal output
rlabel metal3 s 179200 85144 180000 85264 6 b10[21]
port 83 nsew signal output
rlabel metal3 s 0 100104 800 100224 6 b10[22]
port 84 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 b10[23]
port 85 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 b10[24]
port 86 nsew signal output
rlabel metal2 s 122470 119200 122526 120000 6 b10[25]
port 87 nsew signal output
rlabel metal2 s 150898 0 150954 800 6 b10[26]
port 88 nsew signal output
rlabel metal2 s 162030 0 162086 800 6 b10[27]
port 89 nsew signal output
rlabel metal2 s 143078 119200 143134 120000 6 b10[28]
port 90 nsew signal output
rlabel metal3 s 179200 116968 180000 117088 6 b10[29]
port 91 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 b10[2]
port 92 nsew signal output
rlabel metal2 s 170310 0 170366 800 6 b10[30]
port 93 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 b10[31]
port 94 nsew signal output
rlabel metal3 s 179200 17688 180000 17808 6 b10[3]
port 95 nsew signal output
rlabel metal3 s 179200 23264 180000 23384 6 b10[4]
port 96 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 b10[5]
port 97 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 b10[6]
port 98 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 b10[7]
port 99 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 b10[8]
port 100 nsew signal output
rlabel metal3 s 0 52640 800 52760 6 b10[9]
port 101 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 b11[0]
port 102 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 b11[10]
port 103 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 b11[11]
port 104 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 b11[12]
port 105 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 b11[13]
port 106 nsew signal output
rlabel metal3 s 179200 56992 180000 57112 6 b11[14]
port 107 nsew signal output
rlabel metal2 s 81162 119200 81218 120000 6 b11[15]
port 108 nsew signal output
rlabel metal3 s 0 85824 800 85944 6 b11[16]
port 109 nsew signal output
rlabel metal3 s 179200 70048 180000 70168 6 b11[17]
port 110 nsew signal output
rlabel metal3 s 0 87456 800 87576 6 b11[18]
port 111 nsew signal output
rlabel metal3 s 0 90584 800 90704 6 b11[19]
port 112 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 b11[1]
port 113 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 b11[20]
port 114 nsew signal output
rlabel metal3 s 179200 86912 180000 87032 6 b11[21]
port 115 nsew signal output
rlabel metal2 s 107658 119200 107714 120000 6 b11[22]
port 116 nsew signal output
rlabel metal3 s 0 103232 800 103352 6 b11[23]
port 117 nsew signal output
rlabel metal3 s 179200 100104 180000 100224 6 b11[24]
port 118 nsew signal output
rlabel metal2 s 125414 119200 125470 120000 6 b11[25]
port 119 nsew signal output
rlabel metal3 s 179200 109488 180000 109608 6 b11[26]
port 120 nsew signal output
rlabel metal2 s 134246 119200 134302 120000 6 b11[27]
port 121 nsew signal output
rlabel metal2 s 146114 119200 146170 120000 6 b11[28]
port 122 nsew signal output
rlabel metal2 s 157890 119200 157946 120000 6 b11[29]
port 123 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 b11[2]
port 124 nsew signal output
rlabel metal3 s 0 115880 800 116000 6 b11[30]
port 125 nsew signal output
rlabel metal3 s 179200 118872 180000 118992 6 b11[31]
port 126 nsew signal output
rlabel metal2 s 25042 119200 25098 120000 6 b11[3]
port 127 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 b11[4]
port 128 nsew signal output
rlabel metal2 s 39854 119200 39910 120000 6 b11[5]
port 129 nsew signal output
rlabel metal3 s 0 36864 800 36984 6 b11[6]
port 130 nsew signal output
rlabel metal3 s 179200 30744 180000 30864 6 b11[7]
port 131 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 b11[8]
port 132 nsew signal output
rlabel metal3 s 179200 38224 180000 38344 6 b11[9]
port 133 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 b12[0]
port 134 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 b12[10]
port 135 nsew signal output
rlabel metal3 s 0 62160 800 62280 6 b12[11]
port 136 nsew signal output
rlabel metal2 s 72238 119200 72294 120000 6 b12[12]
port 137 nsew signal output
rlabel metal3 s 179200 53184 180000 53304 6 b12[13]
port 138 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 b12[14]
port 139 nsew signal output
rlabel metal2 s 84106 119200 84162 120000 6 b12[15]
port 140 nsew signal output
rlabel metal2 s 89994 119200 90050 120000 6 b12[16]
port 141 nsew signal output
rlabel metal2 s 109406 0 109462 800 6 b12[17]
port 142 nsew signal output
rlabel metal2 s 98826 119200 98882 120000 6 b12[18]
port 143 nsew signal output
rlabel metal3 s 179200 77664 180000 77784 6 b12[19]
port 144 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 b12[1]
port 145 nsew signal output
rlabel metal2 s 137098 0 137154 800 6 b12[20]
port 146 nsew signal output
rlabel metal3 s 179200 88816 180000 88936 6 b12[21]
port 147 nsew signal output
rlabel metal2 s 110694 119200 110750 120000 6 b12[22]
port 148 nsew signal output
rlabel metal2 s 113638 119200 113694 120000 6 b12[23]
port 149 nsew signal output
rlabel metal2 s 145378 0 145434 800 6 b12[24]
port 150 nsew signal output
rlabel metal2 s 128358 119200 128414 120000 6 b12[25]
port 151 nsew signal output
rlabel metal3 s 179200 111392 180000 111512 6 b12[26]
port 152 nsew signal output
rlabel metal2 s 137190 119200 137246 120000 6 b12[27]
port 153 nsew signal output
rlabel metal2 s 149058 119200 149114 120000 6 b12[28]
port 154 nsew signal output
rlabel metal2 s 160834 119200 160890 120000 6 b12[29]
port 155 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 b12[2]
port 156 nsew signal output
rlabel metal3 s 0 117376 800 117496 6 b12[30]
port 157 nsew signal output
rlabel metal2 s 178590 0 178646 800 6 b12[31]
port 158 nsew signal output
rlabel metal2 s 27986 119200 28042 120000 6 b12[3]
port 159 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 b12[4]
port 160 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 b12[5]
port 161 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 b12[6]
port 162 nsew signal output
rlabel metal2 s 54574 119200 54630 120000 6 b12[7]
port 163 nsew signal output
rlabel metal3 s 0 48016 800 48136 6 b12[8]
port 164 nsew signal output
rlabel metal2 s 60462 119200 60518 120000 6 b12[9]
port 165 nsew signal output
rlabel metal3 s 0 688 800 808 6 clk_i
port 166 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 cyc_i
port 167 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 dat_i[0]
port 168 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 dat_i[10]
port 169 nsew signal input
rlabel metal3 s 179200 43800 180000 43920 6 dat_i[11]
port 170 nsew signal input
rlabel metal3 s 0 71680 800 71800 6 dat_i[12]
port 171 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 dat_i[13]
port 172 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 dat_i[14]
port 173 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 dat_i[15]
port 174 nsew signal input
rlabel metal2 s 92938 119200 92994 120000 6 dat_i[16]
port 175 nsew signal input
rlabel metal3 s 179200 71952 180000 72072 6 dat_i[17]
port 176 nsew signal input
rlabel metal3 s 179200 75760 180000 75880 6 dat_i[18]
port 177 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 dat_i[19]
port 178 nsew signal input
rlabel metal2 s 16210 119200 16266 120000 6 dat_i[1]
port 179 nsew signal input
rlabel metal3 s 179200 81336 180000 81456 6 dat_i[20]
port 180 nsew signal input
rlabel metal3 s 179200 90720 180000 90840 6 dat_i[21]
port 181 nsew signal input
rlabel metal3 s 179200 92624 180000 92744 6 dat_i[22]
port 182 nsew signal input
rlabel metal2 s 116582 119200 116638 120000 6 dat_i[23]
port 183 nsew signal input
rlabel metal2 s 119526 119200 119582 120000 6 dat_i[24]
port 184 nsew signal input
rlabel metal3 s 179200 105680 180000 105800 6 dat_i[25]
port 185 nsew signal input
rlabel metal2 s 131302 119200 131358 120000 6 dat_i[26]
port 186 nsew signal input
rlabel metal2 s 164790 0 164846 800 6 dat_i[27]
port 187 nsew signal input
rlabel metal2 s 152002 119200 152058 120000 6 dat_i[28]
port 188 nsew signal input
rlabel metal2 s 163778 119200 163834 120000 6 dat_i[29]
port 189 nsew signal input
rlabel metal3 s 179200 13880 180000 14000 6 dat_i[2]
port 190 nsew signal input
rlabel metal2 s 169666 119200 169722 120000 6 dat_i[30]
port 191 nsew signal input
rlabel metal2 s 175554 119200 175610 120000 6 dat_i[31]
port 192 nsew signal input
rlabel metal2 s 30930 119200 30986 120000 6 dat_i[3]
port 193 nsew signal input
rlabel metal3 s 0 28976 800 29096 6 dat_i[4]
port 194 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 dat_i[5]
port 195 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 dat_i[6]
port 196 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 dat_i[7]
port 197 nsew signal input
rlabel metal3 s 179200 32648 180000 32768 6 dat_i[8]
port 198 nsew signal input
rlabel metal3 s 0 54272 800 54392 6 dat_i[9]
port 199 nsew signal input
rlabel metal2 s 10322 119200 10378 120000 6 dat_o[0]
port 200 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 dat_o[10]
port 201 nsew signal output
rlabel metal3 s 179200 45704 180000 45824 6 dat_o[11]
port 202 nsew signal output
rlabel metal3 s 0 73176 800 73296 6 dat_o[12]
port 203 nsew signal output
rlabel metal3 s 0 76440 800 76560 6 dat_o[13]
port 204 nsew signal output
rlabel metal2 s 95514 0 95570 800 6 dat_o[14]
port 205 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 dat_o[15]
port 206 nsew signal output
rlabel metal3 s 179200 66376 180000 66496 6 dat_o[16]
port 207 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 dat_o[17]
port 208 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 dat_o[18]
port 209 nsew signal output
rlabel metal3 s 179200 79432 180000 79552 6 dat_o[19]
port 210 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 dat_o[1]
port 211 nsew signal output
rlabel metal3 s 0 93712 800 93832 6 dat_o[20]
port 212 nsew signal output
rlabel metal3 s 0 95344 800 95464 6 dat_o[21]
port 213 nsew signal output
rlabel metal3 s 179200 94528 180000 94648 6 dat_o[22]
port 214 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 dat_o[23]
port 215 nsew signal output
rlabel metal3 s 179200 102008 180000 102128 6 dat_o[24]
port 216 nsew signal output
rlabel metal3 s 0 107992 800 108112 6 dat_o[25]
port 217 nsew signal output
rlabel metal2 s 153658 0 153714 800 6 dat_o[26]
port 218 nsew signal output
rlabel metal3 s 0 111120 800 111240 6 dat_o[27]
port 219 nsew signal output
rlabel metal3 s 179200 115064 180000 115184 6 dat_o[28]
port 220 nsew signal output
rlabel metal2 s 166722 119200 166778 120000 6 dat_o[29]
port 221 nsew signal output
rlabel metal2 s 22098 119200 22154 120000 6 dat_o[2]
port 222 nsew signal output
rlabel metal2 s 173070 0 173126 800 6 dat_o[30]
port 223 nsew signal output
rlabel metal2 s 178498 119200 178554 120000 6 dat_o[31]
port 224 nsew signal output
rlabel metal3 s 179200 19456 180000 19576 6 dat_o[3]
port 225 nsew signal output
rlabel metal2 s 36818 119200 36874 120000 6 dat_o[4]
port 226 nsew signal output
rlabel metal2 s 42798 119200 42854 120000 6 dat_o[5]
port 227 nsew signal output
rlabel metal2 s 51630 119200 51686 120000 6 dat_o[6]
port 228 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 dat_o[7]
port 229 nsew signal output
rlabel metal3 s 179200 34552 180000 34672 6 dat_o[8]
port 230 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 dat_o[9]
port 231 nsew signal output
rlabel metal3 s 179200 824 180000 944 6 rst_i
port 232 nsew signal input
rlabel metal3 s 179200 2592 180000 2712 6 stb_i
port 233 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 234 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 234 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 234 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 234 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 234 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 234 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 235 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 235 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 235 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 235 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 235 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 235 nsew ground input
rlabel metal3 s 0 2184 800 2304 6 we_i
port 236 nsew signal input
rlabel metal2 s 13266 119200 13322 120000 6 x[0]
port 237 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 x[10]
port 238 nsew signal input
rlabel metal3 s 0 63792 800 63912 6 x[11]
port 239 nsew signal input
rlabel metal3 s 179200 49512 180000 49632 6 x[12]
port 240 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 x[13]
port 241 nsew signal input
rlabel metal3 s 179200 58896 180000 59016 6 x[14]
port 242 nsew signal input
rlabel metal3 s 0 82696 800 82816 6 x[15]
port 243 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 x[1]
port 244 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 x[2]
port 245 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 x[3]
port 246 nsew signal input
rlabel metal3 s 179200 25168 180000 25288 6 x[4]
port 247 nsew signal input
rlabel metal2 s 45742 119200 45798 120000 6 x[5]
port 248 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 x[6]
port 249 nsew signal input
rlabel metal2 s 57518 119200 57574 120000 6 x[7]
port 250 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 x[8]
port 251 nsew signal input
rlabel metal3 s 0 55904 800 56024 6 x[9]
port 252 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 y[0]
port 253 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 y[10]
port 254 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 y[11]
port 255 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 y[12]
port 256 nsew signal input
rlabel metal3 s 179200 55088 180000 55208 6 y[13]
port 257 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 y[14]
port 258 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 y[15]
port 259 nsew signal input
rlabel metal2 s 19154 119200 19210 120000 6 y[1]
port 260 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 y[2]
port 261 nsew signal input
rlabel metal3 s 179200 21360 180000 21480 6 y[3]
port 262 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 y[4]
port 263 nsew signal input
rlabel metal2 s 48686 119200 48742 120000 6 y[5]
port 264 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 y[6]
port 265 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 y[7]
port 266 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 y[8]
port 267 nsew signal input
rlabel metal3 s 179200 40128 180000 40248 6 y[9]
port 268 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10779592
string GDS_FILE /home/openpdk/caravel/fct-iot-node-project/openlane/coefio/runs/coefio/results/finishing/coefio.magic.gds
string GDS_START 315116
<< end >>

