VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multa
  CLASS BLOCK ;
  FOREIGN multa ;
  ORIGIN 0.000 0.000 ;
  SIZE 272.280 BY 283.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 279.000 168.270 283.000 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 151.000 272.280 151.600 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 191.120 272.280 191.720 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END a[14]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 279.000 8.190 283.000 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 279.000 39.930 283.000 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 279.000 56.030 283.000 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 279.000 88.230 283.000 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 279.000 119.970 283.000 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 70.080 272.280 70.680 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END a[9]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END b[0]
  PIN b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END b[10]
  PIN b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END b[11]
  PIN b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END b[12]
  PIN b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END b[13]
  PIN b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END b[14]
  PIN b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 211.520 272.280 212.120 ;
    END
  END b[15]
  PIN b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END b[16]
  PIN b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 231.240 272.280 231.840 ;
    END
  END b[17]
  PIN b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END b[18]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 9.560 272.280 10.160 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 279.000 72.130 283.000 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 279.000 136.070 283.000 ;
    END
  END b[7]
  PIN b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END b[8]
  PIN b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 110.200 272.280 110.800 ;
    END
  END b[9]
  PIN r[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END r[0]
  PIN r[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END r[10]
  PIN r[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 130.600 272.280 131.200 ;
    END
  END r[11]
  PIN r[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 170.720 272.280 171.320 ;
    END
  END r[12]
  PIN r[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 279.000 184.370 283.000 ;
    END
  END r[13]
  PIN r[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 279.000 200.010 283.000 ;
    END
  END r[14]
  PIN r[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END r[15]
  PIN r[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END r[16]
  PIN r[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END r[17]
  PIN r[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END r[18]
  PIN r[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END r[19]
  PIN r[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END r[1]
  PIN r[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 251.640 272.280 252.240 ;
    END
  END r[20]
  PIN r[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 279.000 216.110 283.000 ;
    END
  END r[21]
  PIN r[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 279.000 232.210 283.000 ;
    END
  END r[22]
  PIN r[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 279.000 248.310 283.000 ;
    END
  END r[23]
  PIN r[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END r[24]
  PIN r[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END r[25]
  PIN r[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END r[26]
  PIN r[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.880 4.000 247.480 ;
    END
  END r[27]
  PIN r[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END r[28]
  PIN r[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END r[29]
  PIN r[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 279.000 23.830 283.000 ;
    END
  END r[2]
  PIN r[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 272.040 272.280 272.640 ;
    END
  END r[30]
  PIN r[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END r[31]
  PIN r[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 279.000 264.410 283.000 ;
    END
  END r[32]
  PIN r[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END r[33]
  PIN r[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 29.280 272.280 29.880 ;
    END
  END r[3]
  PIN r[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END r[4]
  PIN r[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 279.000 103.870 283.000 ;
    END
  END r[5]
  PIN r[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 49.680 272.280 50.280 ;
    END
  END r[6]
  PIN r[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END r[7]
  PIN r[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.280 89.800 272.280 90.400 ;
    END
  END r[8]
  PIN r[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 279.000 152.170 283.000 ;
    END
  END r[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 272.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 272.240 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 266.340 272.085 ;
      LAYER met1 ;
        RECT 5.520 9.560 266.340 272.240 ;
      LAYER met2 ;
        RECT 5.610 278.720 7.630 279.000 ;
        RECT 8.470 278.720 23.270 279.000 ;
        RECT 24.110 278.720 39.370 279.000 ;
        RECT 40.210 278.720 55.470 279.000 ;
        RECT 56.310 278.720 71.570 279.000 ;
        RECT 72.410 278.720 87.670 279.000 ;
        RECT 88.510 278.720 103.310 279.000 ;
        RECT 104.150 278.720 119.410 279.000 ;
        RECT 120.250 278.720 135.510 279.000 ;
        RECT 136.350 278.720 151.610 279.000 ;
        RECT 152.450 278.720 167.710 279.000 ;
        RECT 168.550 278.720 183.810 279.000 ;
        RECT 184.650 278.720 199.450 279.000 ;
        RECT 200.290 278.720 215.550 279.000 ;
        RECT 216.390 278.720 231.650 279.000 ;
        RECT 232.490 278.720 247.750 279.000 ;
        RECT 248.590 278.720 263.850 279.000 ;
        RECT 5.610 4.280 264.400 278.720 ;
        RECT 5.610 4.000 7.630 4.280 ;
        RECT 8.470 4.000 23.270 4.280 ;
        RECT 24.110 4.000 39.370 4.280 ;
        RECT 40.210 4.000 55.470 4.280 ;
        RECT 56.310 4.000 71.570 4.280 ;
        RECT 72.410 4.000 87.670 4.280 ;
        RECT 88.510 4.000 103.310 4.280 ;
        RECT 104.150 4.000 119.410 4.280 ;
        RECT 120.250 4.000 135.510 4.280 ;
        RECT 136.350 4.000 151.610 4.280 ;
        RECT 152.450 4.000 167.710 4.280 ;
        RECT 168.550 4.000 183.810 4.280 ;
        RECT 184.650 4.000 199.450 4.280 ;
        RECT 200.290 4.000 215.550 4.280 ;
        RECT 216.390 4.000 231.650 4.280 ;
        RECT 232.490 4.000 247.750 4.280 ;
        RECT 248.590 4.000 263.850 4.280 ;
      LAYER met3 ;
        RECT 4.400 275.040 268.280 275.905 ;
        RECT 4.000 273.040 268.280 275.040 ;
        RECT 4.000 271.640 267.880 273.040 ;
        RECT 4.000 262.160 268.280 271.640 ;
        RECT 4.400 260.760 268.280 262.160 ;
        RECT 4.000 252.640 268.280 260.760 ;
        RECT 4.000 251.240 267.880 252.640 ;
        RECT 4.000 247.880 268.280 251.240 ;
        RECT 4.400 246.480 268.280 247.880 ;
        RECT 4.000 233.600 268.280 246.480 ;
        RECT 4.400 232.240 268.280 233.600 ;
        RECT 4.400 232.200 267.880 232.240 ;
        RECT 4.000 230.840 267.880 232.200 ;
        RECT 4.000 220.000 268.280 230.840 ;
        RECT 4.400 218.600 268.280 220.000 ;
        RECT 4.000 212.520 268.280 218.600 ;
        RECT 4.000 211.120 267.880 212.520 ;
        RECT 4.000 205.720 268.280 211.120 ;
        RECT 4.400 204.320 268.280 205.720 ;
        RECT 4.000 192.120 268.280 204.320 ;
        RECT 4.000 191.440 267.880 192.120 ;
        RECT 4.400 190.720 267.880 191.440 ;
        RECT 4.400 190.040 268.280 190.720 ;
        RECT 4.000 177.160 268.280 190.040 ;
        RECT 4.400 175.760 268.280 177.160 ;
        RECT 4.000 171.720 268.280 175.760 ;
        RECT 4.000 170.320 267.880 171.720 ;
        RECT 4.000 162.880 268.280 170.320 ;
        RECT 4.400 161.480 268.280 162.880 ;
        RECT 4.000 152.000 268.280 161.480 ;
        RECT 4.000 150.600 267.880 152.000 ;
        RECT 4.000 149.280 268.280 150.600 ;
        RECT 4.400 147.880 268.280 149.280 ;
        RECT 4.000 135.000 268.280 147.880 ;
        RECT 4.400 133.600 268.280 135.000 ;
        RECT 4.000 131.600 268.280 133.600 ;
        RECT 4.000 130.200 267.880 131.600 ;
        RECT 4.000 120.720 268.280 130.200 ;
        RECT 4.400 119.320 268.280 120.720 ;
        RECT 4.000 111.200 268.280 119.320 ;
        RECT 4.000 109.800 267.880 111.200 ;
        RECT 4.000 106.440 268.280 109.800 ;
        RECT 4.400 105.040 268.280 106.440 ;
        RECT 4.000 92.160 268.280 105.040 ;
        RECT 4.400 90.800 268.280 92.160 ;
        RECT 4.400 90.760 267.880 90.800 ;
        RECT 4.000 89.400 267.880 90.760 ;
        RECT 4.000 78.560 268.280 89.400 ;
        RECT 4.400 77.160 268.280 78.560 ;
        RECT 4.000 71.080 268.280 77.160 ;
        RECT 4.000 69.680 267.880 71.080 ;
        RECT 4.000 64.280 268.280 69.680 ;
        RECT 4.400 62.880 268.280 64.280 ;
        RECT 4.000 50.680 268.280 62.880 ;
        RECT 4.000 50.000 267.880 50.680 ;
        RECT 4.400 49.280 267.880 50.000 ;
        RECT 4.400 48.600 268.280 49.280 ;
        RECT 4.000 35.720 268.280 48.600 ;
        RECT 4.400 34.320 268.280 35.720 ;
        RECT 4.000 30.280 268.280 34.320 ;
        RECT 4.000 28.880 267.880 30.280 ;
        RECT 4.000 21.440 268.280 28.880 ;
        RECT 4.400 20.040 268.280 21.440 ;
        RECT 4.000 10.560 268.280 20.040 ;
        RECT 4.000 9.160 267.880 10.560 ;
        RECT 4.000 7.840 268.280 9.160 ;
        RECT 4.400 6.975 268.280 7.840 ;
      LAYER met4 ;
        RECT 12.255 17.175 20.640 269.785 ;
        RECT 23.040 17.175 97.440 269.785 ;
        RECT 99.840 17.175 174.240 269.785 ;
        RECT 176.640 17.175 207.625 269.785 ;
  END
END multa
END LIBRARY

