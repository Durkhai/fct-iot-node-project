magic
tech sky130A
magscale 1 2
timestamp 1653783020
<< obsli1 >>
rect 1104 2159 73692 74545
<< obsm1 >>
rect 1104 1856 73692 74576
<< metal2 >>
rect 2502 76219 2558 77019
rect 7470 76219 7526 77019
rect 12438 76219 12494 77019
rect 17406 76219 17462 77019
rect 22466 76219 22522 77019
rect 27434 76219 27490 77019
rect 32402 76219 32458 77019
rect 37370 76219 37426 77019
rect 42430 76219 42486 77019
rect 47398 76219 47454 77019
rect 52366 76219 52422 77019
rect 57334 76219 57390 77019
rect 62394 76219 62450 77019
rect 67362 76219 67418 77019
rect 72330 76219 72386 77019
rect 2134 0 2190 800
rect 6458 0 6514 800
rect 10874 0 10930 800
rect 15290 0 15346 800
rect 19706 0 19762 800
rect 24122 0 24178 800
rect 28538 0 28594 800
rect 32954 0 33010 800
rect 37370 0 37426 800
rect 41694 0 41750 800
rect 46110 0 46166 800
rect 50526 0 50582 800
rect 54942 0 54998 800
rect 59358 0 59414 800
rect 63774 0 63830 800
rect 68190 0 68246 800
rect 72606 0 72662 800
<< obsm2 >>
rect 1398 76163 2446 76378
rect 2614 76163 7414 76378
rect 7582 76163 12382 76378
rect 12550 76163 17350 76378
rect 17518 76163 22410 76378
rect 22578 76163 27378 76378
rect 27546 76163 32346 76378
rect 32514 76163 37314 76378
rect 37482 76163 42374 76378
rect 42542 76163 47342 76378
rect 47510 76163 52310 76378
rect 52478 76163 57278 76378
rect 57446 76163 62338 76378
rect 62506 76163 67306 76378
rect 67474 76163 72274 76378
rect 72442 76163 73122 76378
rect 1398 856 73122 76163
rect 1398 734 2078 856
rect 2246 734 6402 856
rect 6570 734 10818 856
rect 10986 734 15234 856
rect 15402 734 19650 856
rect 19818 734 24066 856
rect 24234 734 28482 856
rect 28650 734 32898 856
rect 33066 734 37314 856
rect 37482 734 41638 856
rect 41806 734 46054 856
rect 46222 734 50470 856
rect 50638 734 54886 856
rect 55054 734 59302 856
rect 59470 734 63718 856
rect 63886 734 68134 856
rect 68302 734 72550 856
rect 72718 734 73122 856
<< metal3 >>
rect 0 74944 800 75064
rect 74075 75080 74875 75200
rect 74075 71544 74875 71664
rect 0 71136 800 71256
rect 74075 68008 74875 68128
rect 0 67328 800 67448
rect 74075 64608 74875 64728
rect 0 63384 800 63504
rect 74075 61072 74875 61192
rect 0 59576 800 59696
rect 74075 57536 74875 57656
rect 0 55768 800 55888
rect 74075 54000 74875 54120
rect 0 51824 800 51944
rect 74075 50600 74875 50720
rect 0 48016 800 48136
rect 74075 47064 74875 47184
rect 0 44208 800 44328
rect 74075 43528 74875 43648
rect 0 40400 800 40520
rect 74075 40128 74875 40248
rect 0 36456 800 36576
rect 74075 36592 74875 36712
rect 74075 33056 74875 33176
rect 0 32648 800 32768
rect 74075 29520 74875 29640
rect 0 28840 800 28960
rect 74075 26120 74875 26240
rect 0 24896 800 25016
rect 74075 22584 74875 22704
rect 0 21088 800 21208
rect 74075 19048 74875 19168
rect 0 17280 800 17400
rect 74075 15512 74875 15632
rect 0 13336 800 13456
rect 74075 12112 74875 12232
rect 0 9528 800 9648
rect 74075 8576 74875 8696
rect 0 5720 800 5840
rect 74075 5040 74875 5160
rect 0 1912 800 2032
rect 74075 1640 74875 1760
<< obsm3 >>
rect 800 75144 73995 75173
rect 880 75000 73995 75144
rect 880 74864 74075 75000
rect 800 71744 74075 74864
rect 800 71464 73995 71744
rect 800 71336 74075 71464
rect 880 71056 74075 71336
rect 800 68208 74075 71056
rect 800 67928 73995 68208
rect 800 67528 74075 67928
rect 880 67248 74075 67528
rect 800 64808 74075 67248
rect 800 64528 73995 64808
rect 800 63584 74075 64528
rect 880 63304 74075 63584
rect 800 61272 74075 63304
rect 800 60992 73995 61272
rect 800 59776 74075 60992
rect 880 59496 74075 59776
rect 800 57736 74075 59496
rect 800 57456 73995 57736
rect 800 55968 74075 57456
rect 880 55688 74075 55968
rect 800 54200 74075 55688
rect 800 53920 73995 54200
rect 800 52024 74075 53920
rect 880 51744 74075 52024
rect 800 50800 74075 51744
rect 800 50520 73995 50800
rect 800 48216 74075 50520
rect 880 47936 74075 48216
rect 800 47264 74075 47936
rect 800 46984 73995 47264
rect 800 44408 74075 46984
rect 880 44128 74075 44408
rect 800 43728 74075 44128
rect 800 43448 73995 43728
rect 800 40600 74075 43448
rect 880 40328 74075 40600
rect 880 40320 73995 40328
rect 800 40048 73995 40320
rect 800 36792 74075 40048
rect 800 36656 73995 36792
rect 880 36512 73995 36656
rect 880 36376 74075 36512
rect 800 33256 74075 36376
rect 800 32976 73995 33256
rect 800 32848 74075 32976
rect 880 32568 74075 32848
rect 800 29720 74075 32568
rect 800 29440 73995 29720
rect 800 29040 74075 29440
rect 880 28760 74075 29040
rect 800 26320 74075 28760
rect 800 26040 73995 26320
rect 800 25096 74075 26040
rect 880 24816 74075 25096
rect 800 22784 74075 24816
rect 800 22504 73995 22784
rect 800 21288 74075 22504
rect 880 21008 74075 21288
rect 800 19248 74075 21008
rect 800 18968 73995 19248
rect 800 17480 74075 18968
rect 880 17200 74075 17480
rect 800 15712 74075 17200
rect 800 15432 73995 15712
rect 800 13536 74075 15432
rect 880 13256 74075 13536
rect 800 12312 74075 13256
rect 800 12032 73995 12312
rect 800 9728 74075 12032
rect 880 9448 74075 9728
rect 800 8776 74075 9448
rect 800 8496 73995 8776
rect 800 5920 74075 8496
rect 880 5640 74075 5920
rect 800 5240 74075 5640
rect 800 4960 73995 5240
rect 800 2112 74075 4960
rect 880 1840 74075 2112
rect 880 1832 73995 1840
rect 800 1667 73995 1832
<< metal4 >>
rect 4208 2128 4528 74576
rect 19568 2128 19888 74576
rect 34928 2128 35248 74576
rect 50288 2128 50608 74576
rect 65648 2128 65968 74576
<< obsm4 >>
rect 9443 2347 19488 74221
rect 19968 2347 34848 74221
rect 35328 2347 50208 74221
rect 50688 2347 65568 74221
rect 66048 2347 72805 74221
<< labels >>
rlabel metal2 s 6458 0 6514 800 6 a11[0]
port 1 nsew signal input
rlabel metal3 s 74075 5040 74875 5160 6 a11[1]
port 2 nsew signal input
rlabel metal3 s 74075 12112 74875 12232 6 a11[2]
port 3 nsew signal input
rlabel metal2 s 22466 76219 22522 77019 6 a11[3]
port 4 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 a11[4]
port 5 nsew signal input
rlabel metal3 s 74075 36592 74875 36712 6 a11[5]
port 6 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 a11[6]
port 7 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 a11[7]
port 8 nsew signal input
rlabel metal3 s 0 71136 800 71256 6 a11[8]
port 9 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 a11[9]
port 10 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 a12[0]
port 11 nsew signal input
rlabel metal2 s 7470 76219 7526 77019 6 a12[1]
port 12 nsew signal input
rlabel metal3 s 74075 15512 74875 15632 6 a12[2]
port 13 nsew signal input
rlabel metal2 s 27434 76219 27490 77019 6 a12[3]
port 14 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 a12[4]
port 15 nsew signal input
rlabel metal3 s 74075 40128 74875 40248 6 a12[5]
port 16 nsew signal input
rlabel metal3 s 74075 47064 74875 47184 6 a12[6]
port 17 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 a12[7]
port 18 nsew signal input
rlabel metal2 s 57334 76219 57390 77019 6 a12[8]
port 19 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 a12[9]
port 20 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 b10[0]
port 21 nsew signal input
rlabel metal2 s 12438 76219 12494 77019 6 b10[1]
port 22 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 b10[2]
port 23 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 b10[3]
port 24 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 b10[4]
port 25 nsew signal input
rlabel metal3 s 0 48016 800 48136 6 b10[5]
port 26 nsew signal input
rlabel metal2 s 47398 76219 47454 77019 6 b10[6]
port 27 nsew signal input
rlabel metal3 s 74075 57536 74875 57656 6 b10[7]
port 28 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 b10[8]
port 29 nsew signal input
rlabel metal3 s 74075 71544 74875 71664 6 b10[9]
port 30 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 b11[0]
port 31 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 b11[1]
port 32 nsew signal input
rlabel metal3 s 74075 19048 74875 19168 6 b11[2]
port 33 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 b11[3]
port 34 nsew signal input
rlabel metal3 s 74075 29520 74875 29640 6 b11[4]
port 35 nsew signal input
rlabel metal2 s 37370 76219 37426 77019 6 b11[5]
port 36 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 b11[6]
port 37 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 b11[7]
port 38 nsew signal input
rlabel metal2 s 62394 76219 62450 77019 6 b11[8]
port 39 nsew signal input
rlabel metal3 s 74075 75080 74875 75200 6 b11[9]
port 40 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 b12[0]
port 41 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 b12[1]
port 42 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 b12[2]
port 43 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 b12[3]
port 44 nsew signal input
rlabel metal3 s 74075 33056 74875 33176 6 b12[4]
port 45 nsew signal input
rlabel metal2 s 42430 76219 42486 77019 6 b12[5]
port 46 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 b12[6]
port 47 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 b12[7]
port 48 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 b12[8]
port 49 nsew signal input
rlabel metal2 s 67362 76219 67418 77019 6 b12[9]
port 50 nsew signal input
rlabel metal2 s 2502 76219 2558 77019 6 clk
port 51 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 enable
port 52 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 nreset
port 53 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 valid
port 54 nsew signal input
rlabel metal4 s 4208 2128 4528 74576 6 vccd1
port 55 nsew power input
rlabel metal4 s 34928 2128 35248 74576 6 vccd1
port 55 nsew power input
rlabel metal4 s 65648 2128 65968 74576 6 vccd1
port 55 nsew power input
rlabel metal4 s 19568 2128 19888 74576 6 vssd1
port 56 nsew ground input
rlabel metal4 s 50288 2128 50608 74576 6 vssd1
port 56 nsew ground input
rlabel metal3 s 0 17280 800 17400 6 x[0]
port 57 nsew signal input
rlabel metal2 s 17406 76219 17462 77019 6 x[1]
port 58 nsew signal input
rlabel metal3 s 74075 22584 74875 22704 6 x[2]
port 59 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 x[3]
port 60 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 x[4]
port 61 nsew signal input
rlabel metal3 s 74075 43528 74875 43648 6 x[5]
port 62 nsew signal input
rlabel metal3 s 74075 50600 74875 50720 6 x[6]
port 63 nsew signal input
rlabel metal3 s 74075 61072 74875 61192 6 x[7]
port 64 nsew signal input
rlabel metal3 s 74075 64608 74875 64728 6 x[8]
port 65 nsew signal input
rlabel metal2 s 72330 76219 72386 77019 6 x[9]
port 66 nsew signal input
rlabel metal3 s 74075 1640 74875 1760 6 yout[0]
port 67 nsew signal output
rlabel metal3 s 74075 8576 74875 8696 6 yout[1]
port 68 nsew signal output
rlabel metal3 s 74075 26120 74875 26240 6 yout[2]
port 69 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 yout[3]
port 70 nsew signal output
rlabel metal2 s 32402 76219 32458 77019 6 yout[4]
port 71 nsew signal output
rlabel metal3 s 0 51824 800 51944 6 yout[5]
port 72 nsew signal output
rlabel metal3 s 74075 54000 74875 54120 6 yout[6]
port 73 nsew signal output
rlabel metal2 s 52366 76219 52422 77019 6 yout[7]
port 74 nsew signal output
rlabel metal3 s 74075 68008 74875 68128 6 yout[8]
port 75 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 yout[9]
port 76 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 74875 77019
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 14673958
string GDS_FILE /home/openpdk/caravel/fct-iot-node-project/openlane/biquad/runs/biquad/results/finishing/biquad.magic.gds
string GDS_START 755186
<< end >>

