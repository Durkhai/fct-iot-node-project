magic
tech sky130A
magscale 1 2
timestamp 1654717483
<< nwell >>
rect 1066 212421 282202 212742
rect 1066 211333 282202 211899
rect 1066 210245 282202 210811
rect 1066 209157 282202 209723
rect 1066 208069 282202 208635
rect 1066 206981 282202 207547
rect 1066 205893 282202 206459
rect 1066 204805 282202 205371
rect 1066 203717 282202 204283
rect 1066 202629 282202 203195
rect 1066 201541 282202 202107
rect 1066 200453 282202 201019
rect 1066 199365 282202 199931
rect 1066 198277 282202 198843
rect 1066 197189 282202 197755
rect 1066 196101 282202 196667
rect 1066 195013 282202 195579
rect 1066 193925 282202 194491
rect 1066 192837 282202 193403
rect 1066 191749 282202 192315
rect 1066 190661 282202 191227
rect 1066 189573 282202 190139
rect 1066 188485 282202 189051
rect 1066 187397 282202 187963
rect 1066 186309 282202 186875
rect 1066 185221 282202 185787
rect 1066 184133 282202 184699
rect 1066 183045 282202 183611
rect 1066 181957 282202 182523
rect 1066 180869 282202 181435
rect 1066 179781 282202 180347
rect 1066 178693 282202 179259
rect 1066 177605 282202 178171
rect 1066 176517 282202 177083
rect 1066 175429 282202 175995
rect 1066 174341 282202 174907
rect 1066 173253 282202 173819
rect 1066 172165 282202 172731
rect 1066 171077 282202 171643
rect 1066 169989 282202 170555
rect 1066 168901 282202 169467
rect 1066 167813 282202 168379
rect 1066 166725 282202 167291
rect 1066 165637 282202 166203
rect 1066 164549 282202 165115
rect 1066 163461 282202 164027
rect 1066 162373 282202 162939
rect 1066 161285 282202 161851
rect 1066 160197 282202 160763
rect 1066 159109 282202 159675
rect 1066 158021 282202 158587
rect 1066 156933 282202 157499
rect 1066 155845 282202 156411
rect 1066 154757 282202 155323
rect 1066 153669 282202 154235
rect 1066 152581 282202 153147
rect 1066 151493 282202 152059
rect 1066 150405 282202 150971
rect 1066 149317 282202 149883
rect 1066 148229 282202 148795
rect 1066 147141 282202 147707
rect 1066 146053 282202 146619
rect 1066 144965 282202 145531
rect 1066 143877 282202 144443
rect 1066 142789 282202 143355
rect 1066 141701 282202 142267
rect 1066 140613 282202 141179
rect 1066 139525 282202 140091
rect 1066 138437 282202 139003
rect 1066 137349 282202 137915
rect 1066 136261 282202 136827
rect 1066 135173 282202 135739
rect 1066 134085 282202 134651
rect 1066 132997 282202 133563
rect 1066 131909 282202 132475
rect 1066 130821 282202 131387
rect 1066 129733 282202 130299
rect 1066 128645 282202 129211
rect 1066 127557 282202 128123
rect 1066 126469 282202 127035
rect 1066 125381 282202 125947
rect 1066 124293 282202 124859
rect 1066 123205 282202 123771
rect 1066 122117 282202 122683
rect 1066 121029 282202 121595
rect 1066 119941 282202 120507
rect 1066 118853 282202 119419
rect 1066 117765 282202 118331
rect 1066 116677 282202 117243
rect 1066 115589 282202 116155
rect 1066 114501 282202 115067
rect 1066 113413 282202 113979
rect 1066 112325 282202 112891
rect 1066 111237 282202 111803
rect 1066 110149 282202 110715
rect 1066 109061 282202 109627
rect 1066 107973 282202 108539
rect 1066 106885 282202 107451
rect 1066 105797 282202 106363
rect 1066 104709 282202 105275
rect 1066 103621 282202 104187
rect 1066 102533 282202 103099
rect 1066 101445 282202 102011
rect 1066 100357 282202 100923
rect 1066 99269 282202 99835
rect 1066 98181 282202 98747
rect 1066 97093 282202 97659
rect 1066 96005 282202 96571
rect 1066 94917 282202 95483
rect 1066 93829 282202 94395
rect 1066 92741 282202 93307
rect 1066 91653 282202 92219
rect 1066 90565 282202 91131
rect 1066 89477 282202 90043
rect 1066 88389 282202 88955
rect 1066 87301 282202 87867
rect 1066 86213 282202 86779
rect 1066 85125 282202 85691
rect 1066 84037 282202 84603
rect 1066 82949 282202 83515
rect 1066 81861 282202 82427
rect 1066 80773 282202 81339
rect 1066 79685 282202 80251
rect 1066 78597 282202 79163
rect 1066 77509 282202 78075
rect 1066 76421 282202 76987
rect 1066 75333 282202 75899
rect 1066 74245 282202 74811
rect 1066 73157 282202 73723
rect 1066 72069 282202 72635
rect 1066 70981 282202 71547
rect 1066 69893 282202 70459
rect 1066 68805 282202 69371
rect 1066 67717 282202 68283
rect 1066 66629 282202 67195
rect 1066 65541 282202 66107
rect 1066 64453 282202 65019
rect 1066 63365 282202 63931
rect 1066 62277 282202 62843
rect 1066 61189 282202 61755
rect 1066 60101 282202 60667
rect 1066 59013 282202 59579
rect 1066 57925 282202 58491
rect 1066 56837 282202 57403
rect 1066 55749 282202 56315
rect 1066 54661 282202 55227
rect 1066 53573 282202 54139
rect 1066 52485 282202 53051
rect 1066 51397 282202 51963
rect 1066 50309 282202 50875
rect 1066 49221 282202 49787
rect 1066 48133 282202 48699
rect 1066 47045 282202 47611
rect 1066 45957 282202 46523
rect 1066 44869 282202 45435
rect 1066 43781 282202 44347
rect 1066 42693 282202 43259
rect 1066 41605 282202 42171
rect 1066 40517 282202 41083
rect 1066 39429 282202 39995
rect 1066 38341 282202 38907
rect 1066 37253 282202 37819
rect 1066 36165 282202 36731
rect 1066 35077 282202 35643
rect 1066 33989 282202 34555
rect 1066 32901 282202 33467
rect 1066 31813 282202 32379
rect 1066 30725 282202 31291
rect 1066 29637 282202 30203
rect 1066 28549 282202 29115
rect 1066 27461 282202 28027
rect 1066 26373 282202 26939
rect 1066 25285 282202 25851
rect 1066 24197 282202 24763
rect 1066 23109 282202 23675
rect 1066 22021 282202 22587
rect 1066 20933 282202 21499
rect 1066 19845 282202 20411
rect 1066 18757 282202 19323
rect 1066 17669 282202 18235
rect 1066 16581 282202 17147
rect 1066 15493 282202 16059
rect 1066 14405 282202 14971
rect 1066 13317 282202 13883
rect 1066 12229 282202 12795
rect 1066 11141 282202 11707
rect 1066 10053 282202 10619
rect 1066 8965 282202 9531
rect 1066 7877 282202 8443
rect 1066 6789 282202 7355
rect 1066 5701 282202 6267
rect 1066 4613 282202 5179
rect 1066 3525 282202 4091
rect 1066 2437 282202 3003
<< obsli1 >>
rect 1104 2159 282164 212721
<< obsm1 >>
rect 1104 1776 282164 212752
<< metal2 >>
rect 7838 214390 7894 215190
rect 23570 214390 23626 215190
rect 39302 214390 39358 215190
rect 55034 214390 55090 215190
rect 70766 214390 70822 215190
rect 86498 214390 86554 215190
rect 102230 214390 102286 215190
rect 117962 214390 118018 215190
rect 133694 214390 133750 215190
rect 149518 214390 149574 215190
rect 165250 214390 165306 215190
rect 180982 214390 181038 215190
rect 196714 214390 196770 215190
rect 212446 214390 212502 215190
rect 228178 214390 228234 215190
rect 243910 214390 243966 215190
rect 259642 214390 259698 215190
rect 275374 214390 275430 215190
rect 1306 0 1362 800
rect 3974 0 4030 800
rect 6734 0 6790 800
rect 9494 0 9550 800
rect 12254 0 12310 800
rect 15014 0 15070 800
rect 17774 0 17830 800
rect 20534 0 20590 800
rect 23294 0 23350 800
rect 26054 0 26110 800
rect 28814 0 28870 800
rect 31482 0 31538 800
rect 34242 0 34298 800
rect 37002 0 37058 800
rect 39762 0 39818 800
rect 42522 0 42578 800
rect 45282 0 45338 800
rect 48042 0 48098 800
rect 50802 0 50858 800
rect 53562 0 53618 800
rect 56322 0 56378 800
rect 58990 0 59046 800
rect 61750 0 61806 800
rect 64510 0 64566 800
rect 67270 0 67326 800
rect 70030 0 70086 800
rect 72790 0 72846 800
rect 75550 0 75606 800
rect 78310 0 78366 800
rect 81070 0 81126 800
rect 83830 0 83886 800
rect 86498 0 86554 800
rect 89258 0 89314 800
rect 92018 0 92074 800
rect 94778 0 94834 800
rect 97538 0 97594 800
rect 100298 0 100354 800
rect 103058 0 103114 800
rect 105818 0 105874 800
rect 108578 0 108634 800
rect 111338 0 111394 800
rect 114098 0 114154 800
rect 116766 0 116822 800
rect 119526 0 119582 800
rect 122286 0 122342 800
rect 125046 0 125102 800
rect 127806 0 127862 800
rect 130566 0 130622 800
rect 133326 0 133382 800
rect 136086 0 136142 800
rect 138846 0 138902 800
rect 141606 0 141662 800
rect 144274 0 144330 800
rect 147034 0 147090 800
rect 149794 0 149850 800
rect 152554 0 152610 800
rect 155314 0 155370 800
rect 158074 0 158130 800
rect 160834 0 160890 800
rect 163594 0 163650 800
rect 166354 0 166410 800
rect 169114 0 169170 800
rect 171782 0 171838 800
rect 174542 0 174598 800
rect 177302 0 177358 800
rect 180062 0 180118 800
rect 182822 0 182878 800
rect 185582 0 185638 800
rect 188342 0 188398 800
rect 191102 0 191158 800
rect 193862 0 193918 800
rect 196622 0 196678 800
rect 199382 0 199438 800
rect 202050 0 202106 800
rect 204810 0 204866 800
rect 207570 0 207626 800
rect 210330 0 210386 800
rect 213090 0 213146 800
rect 215850 0 215906 800
rect 218610 0 218666 800
rect 221370 0 221426 800
rect 224130 0 224186 800
rect 226890 0 226946 800
rect 229558 0 229614 800
rect 232318 0 232374 800
rect 235078 0 235134 800
rect 237838 0 237894 800
rect 240598 0 240654 800
rect 243358 0 243414 800
rect 246118 0 246174 800
rect 248878 0 248934 800
rect 251638 0 251694 800
rect 254398 0 254454 800
rect 257066 0 257122 800
rect 259826 0 259882 800
rect 262586 0 262642 800
rect 265346 0 265402 800
rect 268106 0 268162 800
rect 270866 0 270922 800
rect 273626 0 273682 800
rect 276386 0 276442 800
rect 279146 0 279202 800
rect 281906 0 281962 800
<< obsm2 >>
rect 1308 214334 7782 214418
rect 7950 214334 23514 214418
rect 23682 214334 39246 214418
rect 39414 214334 54978 214418
rect 55146 214334 70710 214418
rect 70878 214334 86442 214418
rect 86610 214334 102174 214418
rect 102342 214334 117906 214418
rect 118074 214334 133638 214418
rect 133806 214334 149462 214418
rect 149630 214334 165194 214418
rect 165362 214334 180926 214418
rect 181094 214334 196658 214418
rect 196826 214334 212390 214418
rect 212558 214334 228122 214418
rect 228290 214334 243854 214418
rect 244022 214334 259586 214418
rect 259754 214334 275318 214418
rect 275486 214334 281960 214418
rect 1308 856 281960 214334
rect 1418 734 3918 856
rect 4086 734 6678 856
rect 6846 734 9438 856
rect 9606 734 12198 856
rect 12366 734 14958 856
rect 15126 734 17718 856
rect 17886 734 20478 856
rect 20646 734 23238 856
rect 23406 734 25998 856
rect 26166 734 28758 856
rect 28926 734 31426 856
rect 31594 734 34186 856
rect 34354 734 36946 856
rect 37114 734 39706 856
rect 39874 734 42466 856
rect 42634 734 45226 856
rect 45394 734 47986 856
rect 48154 734 50746 856
rect 50914 734 53506 856
rect 53674 734 56266 856
rect 56434 734 58934 856
rect 59102 734 61694 856
rect 61862 734 64454 856
rect 64622 734 67214 856
rect 67382 734 69974 856
rect 70142 734 72734 856
rect 72902 734 75494 856
rect 75662 734 78254 856
rect 78422 734 81014 856
rect 81182 734 83774 856
rect 83942 734 86442 856
rect 86610 734 89202 856
rect 89370 734 91962 856
rect 92130 734 94722 856
rect 94890 734 97482 856
rect 97650 734 100242 856
rect 100410 734 103002 856
rect 103170 734 105762 856
rect 105930 734 108522 856
rect 108690 734 111282 856
rect 111450 734 114042 856
rect 114210 734 116710 856
rect 116878 734 119470 856
rect 119638 734 122230 856
rect 122398 734 124990 856
rect 125158 734 127750 856
rect 127918 734 130510 856
rect 130678 734 133270 856
rect 133438 734 136030 856
rect 136198 734 138790 856
rect 138958 734 141550 856
rect 141718 734 144218 856
rect 144386 734 146978 856
rect 147146 734 149738 856
rect 149906 734 152498 856
rect 152666 734 155258 856
rect 155426 734 158018 856
rect 158186 734 160778 856
rect 160946 734 163538 856
rect 163706 734 166298 856
rect 166466 734 169058 856
rect 169226 734 171726 856
rect 171894 734 174486 856
rect 174654 734 177246 856
rect 177414 734 180006 856
rect 180174 734 182766 856
rect 182934 734 185526 856
rect 185694 734 188286 856
rect 188454 734 191046 856
rect 191214 734 193806 856
rect 193974 734 196566 856
rect 196734 734 199326 856
rect 199494 734 201994 856
rect 202162 734 204754 856
rect 204922 734 207514 856
rect 207682 734 210274 856
rect 210442 734 213034 856
rect 213202 734 215794 856
rect 215962 734 218554 856
rect 218722 734 221314 856
rect 221482 734 224074 856
rect 224242 734 226834 856
rect 227002 734 229502 856
rect 229670 734 232262 856
rect 232430 734 235022 856
rect 235190 734 237782 856
rect 237950 734 240542 856
rect 240710 734 243302 856
rect 243470 734 246062 856
rect 246230 734 248822 856
rect 248990 734 251582 856
rect 251750 734 254342 856
rect 254510 734 257010 856
rect 257178 734 259770 856
rect 259938 734 262530 856
rect 262698 734 265290 856
rect 265458 734 268050 856
rect 268218 734 270810 856
rect 270978 734 273570 856
rect 273738 734 276330 856
rect 276498 734 279090 856
rect 279258 734 281850 856
<< metal3 >>
rect 282526 208360 283326 208480
rect 282526 194896 283326 195016
rect 282526 181432 283326 181552
rect 282526 167968 283326 168088
rect 282526 154504 283326 154624
rect 282526 141040 283326 141160
rect 282526 127576 283326 127696
rect 282526 114248 283326 114368
rect 282526 100784 283326 100904
rect 282526 87320 283326 87440
rect 282526 73856 283326 73976
rect 282526 60392 283326 60512
rect 282526 46928 283326 47048
rect 282526 33464 283326 33584
rect 282526 20000 283326 20120
rect 282526 6672 283326 6792
<< obsm3 >>
rect 4208 208560 282526 212737
rect 4208 208280 282446 208560
rect 4208 195096 282526 208280
rect 4208 194816 282446 195096
rect 4208 181632 282526 194816
rect 4208 181352 282446 181632
rect 4208 168168 282526 181352
rect 4208 167888 282446 168168
rect 4208 154704 282526 167888
rect 4208 154424 282446 154704
rect 4208 141240 282526 154424
rect 4208 140960 282446 141240
rect 4208 127776 282526 140960
rect 4208 127496 282446 127776
rect 4208 114448 282526 127496
rect 4208 114168 282446 114448
rect 4208 100984 282526 114168
rect 4208 100704 282446 100984
rect 4208 87520 282526 100704
rect 4208 87240 282446 87520
rect 4208 74056 282526 87240
rect 4208 73776 282446 74056
rect 4208 60592 282526 73776
rect 4208 60312 282446 60592
rect 4208 47128 282526 60312
rect 4208 46848 282446 47128
rect 4208 33664 282526 46848
rect 4208 33384 282446 33664
rect 4208 20200 282526 33384
rect 4208 19920 282446 20200
rect 4208 6872 282526 19920
rect 4208 6592 282446 6872
rect 4208 2143 282526 6592
<< metal4 >>
rect 4208 2128 4528 212752
rect 19568 2128 19888 212752
rect 34928 2128 35248 212752
rect 50288 2128 50608 212752
rect 65648 2128 65968 212752
rect 81008 2128 81328 212752
rect 96368 2128 96688 212752
rect 111728 2128 112048 212752
rect 127088 2128 127408 212752
rect 142448 2128 142768 212752
rect 157808 2128 158128 212752
rect 173168 2128 173488 212752
rect 188528 2128 188848 212752
rect 203888 2128 204208 212752
rect 219248 2128 219568 212752
rect 234608 2128 234928 212752
rect 249968 2128 250288 212752
rect 265328 2128 265648 212752
rect 280688 2128 281008 212752
<< obsm4 >>
rect 38331 8875 50208 212397
rect 50688 8875 65568 212397
rect 66048 8875 80928 212397
rect 81408 8875 96288 212397
rect 96768 8875 111648 212397
rect 112128 8875 127008 212397
rect 127488 8875 142368 212397
rect 142848 8875 157728 212397
rect 158208 8875 173088 212397
rect 173568 8875 188448 212397
rect 188928 8875 203808 212397
rect 204288 8875 219168 212397
rect 219648 8875 234528 212397
rect 235008 8875 249888 212397
rect 250368 8875 250549 212397
<< labels >>
rlabel metal2 s 281906 0 281962 800 6 bq_clk_i
port 1 nsew signal input
rlabel metal2 s 7838 214390 7894 215190 6 nreset
port 2 nsew signal input
rlabel metal2 s 23570 214390 23626 215190 6 valid_i
port 3 nsew signal input
rlabel metal4 s 4208 2128 4528 212752 6 vccd1
port 4 nsew power input
rlabel metal4 s 34928 2128 35248 212752 6 vccd1
port 4 nsew power input
rlabel metal4 s 65648 2128 65968 212752 6 vccd1
port 4 nsew power input
rlabel metal4 s 96368 2128 96688 212752 6 vccd1
port 4 nsew power input
rlabel metal4 s 127088 2128 127408 212752 6 vccd1
port 4 nsew power input
rlabel metal4 s 157808 2128 158128 212752 6 vccd1
port 4 nsew power input
rlabel metal4 s 188528 2128 188848 212752 6 vccd1
port 4 nsew power input
rlabel metal4 s 219248 2128 219568 212752 6 vccd1
port 4 nsew power input
rlabel metal4 s 249968 2128 250288 212752 6 vccd1
port 4 nsew power input
rlabel metal4 s 280688 2128 281008 212752 6 vccd1
port 4 nsew power input
rlabel metal4 s 19568 2128 19888 212752 6 vssd1
port 5 nsew ground input
rlabel metal4 s 50288 2128 50608 212752 6 vssd1
port 5 nsew ground input
rlabel metal4 s 81008 2128 81328 212752 6 vssd1
port 5 nsew ground input
rlabel metal4 s 111728 2128 112048 212752 6 vssd1
port 5 nsew ground input
rlabel metal4 s 142448 2128 142768 212752 6 vssd1
port 5 nsew ground input
rlabel metal4 s 173168 2128 173488 212752 6 vssd1
port 5 nsew ground input
rlabel metal4 s 203888 2128 204208 212752 6 vssd1
port 5 nsew ground input
rlabel metal4 s 234608 2128 234928 212752 6 vssd1
port 5 nsew ground input
rlabel metal4 s 265328 2128 265648 212752 6 vssd1
port 5 nsew ground input
rlabel metal2 s 1306 0 1362 800 6 wb_ack_o
port 6 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wb_adr_i[0]
port 7 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 wb_adr_i[10]
port 8 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 wb_adr_i[11]
port 9 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 wb_adr_i[12]
port 10 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 wb_adr_i[13]
port 11 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 wb_adr_i[14]
port 12 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 wb_adr_i[15]
port 13 nsew signal input
rlabel metal2 s 149794 0 149850 800 6 wb_adr_i[16]
port 14 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 wb_adr_i[17]
port 15 nsew signal input
rlabel metal2 s 166354 0 166410 800 6 wb_adr_i[18]
port 16 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 wb_adr_i[19]
port 17 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wb_adr_i[1]
port 18 nsew signal input
rlabel metal2 s 182822 0 182878 800 6 wb_adr_i[20]
port 19 nsew signal input
rlabel metal2 s 191102 0 191158 800 6 wb_adr_i[21]
port 20 nsew signal input
rlabel metal2 s 199382 0 199438 800 6 wb_adr_i[22]
port 21 nsew signal input
rlabel metal2 s 207570 0 207626 800 6 wb_adr_i[23]
port 22 nsew signal input
rlabel metal2 s 215850 0 215906 800 6 wb_adr_i[24]
port 23 nsew signal input
rlabel metal2 s 224130 0 224186 800 6 wb_adr_i[25]
port 24 nsew signal input
rlabel metal2 s 232318 0 232374 800 6 wb_adr_i[26]
port 25 nsew signal input
rlabel metal2 s 240598 0 240654 800 6 wb_adr_i[27]
port 26 nsew signal input
rlabel metal2 s 248878 0 248934 800 6 wb_adr_i[28]
port 27 nsew signal input
rlabel metal2 s 257066 0 257122 800 6 wb_adr_i[29]
port 28 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wb_adr_i[2]
port 29 nsew signal input
rlabel metal2 s 265346 0 265402 800 6 wb_adr_i[30]
port 30 nsew signal input
rlabel metal2 s 273626 0 273682 800 6 wb_adr_i[31]
port 31 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wb_adr_i[3]
port 32 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wb_adr_i[4]
port 33 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 wb_adr_i[5]
port 34 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 wb_adr_i[6]
port 35 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 wb_adr_i[7]
port 36 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 wb_adr_i[8]
port 37 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 wb_adr_i[9]
port 38 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wb_clk_i
port 39 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wb_cyc_i
port 40 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wb_dat_i[0]
port 41 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 wb_dat_i[10]
port 42 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 wb_dat_i[11]
port 43 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 wb_dat_i[12]
port 44 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 wb_dat_i[13]
port 45 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 wb_dat_i[14]
port 46 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 wb_dat_i[15]
port 47 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 wb_dat_i[16]
port 48 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 wb_dat_i[17]
port 49 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 wb_dat_i[18]
port 50 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 wb_dat_i[19]
port 51 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wb_dat_i[1]
port 52 nsew signal input
rlabel metal2 s 185582 0 185638 800 6 wb_dat_i[20]
port 53 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 wb_dat_i[21]
port 54 nsew signal input
rlabel metal2 s 202050 0 202106 800 6 wb_dat_i[22]
port 55 nsew signal input
rlabel metal2 s 210330 0 210386 800 6 wb_dat_i[23]
port 56 nsew signal input
rlabel metal2 s 218610 0 218666 800 6 wb_dat_i[24]
port 57 nsew signal input
rlabel metal2 s 226890 0 226946 800 6 wb_dat_i[25]
port 58 nsew signal input
rlabel metal2 s 235078 0 235134 800 6 wb_dat_i[26]
port 59 nsew signal input
rlabel metal2 s 243358 0 243414 800 6 wb_dat_i[27]
port 60 nsew signal input
rlabel metal2 s 251638 0 251694 800 6 wb_dat_i[28]
port 61 nsew signal input
rlabel metal2 s 259826 0 259882 800 6 wb_dat_i[29]
port 62 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wb_dat_i[2]
port 63 nsew signal input
rlabel metal2 s 268106 0 268162 800 6 wb_dat_i[30]
port 64 nsew signal input
rlabel metal2 s 276386 0 276442 800 6 wb_dat_i[31]
port 65 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wb_dat_i[3]
port 66 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 wb_dat_i[4]
port 67 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 wb_dat_i[5]
port 68 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 wb_dat_i[6]
port 69 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 wb_dat_i[7]
port 70 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 wb_dat_i[8]
port 71 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 wb_dat_i[9]
port 72 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wb_dat_o[0]
port 73 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 wb_dat_o[10]
port 74 nsew signal output
rlabel metal2 s 114098 0 114154 800 6 wb_dat_o[11]
port 75 nsew signal output
rlabel metal2 s 122286 0 122342 800 6 wb_dat_o[12]
port 76 nsew signal output
rlabel metal2 s 130566 0 130622 800 6 wb_dat_o[13]
port 77 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 wb_dat_o[14]
port 78 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 wb_dat_o[15]
port 79 nsew signal output
rlabel metal2 s 155314 0 155370 800 6 wb_dat_o[16]
port 80 nsew signal output
rlabel metal2 s 163594 0 163650 800 6 wb_dat_o[17]
port 81 nsew signal output
rlabel metal2 s 171782 0 171838 800 6 wb_dat_o[18]
port 82 nsew signal output
rlabel metal2 s 180062 0 180118 800 6 wb_dat_o[19]
port 83 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 wb_dat_o[1]
port 84 nsew signal output
rlabel metal2 s 188342 0 188398 800 6 wb_dat_o[20]
port 85 nsew signal output
rlabel metal2 s 196622 0 196678 800 6 wb_dat_o[21]
port 86 nsew signal output
rlabel metal2 s 204810 0 204866 800 6 wb_dat_o[22]
port 87 nsew signal output
rlabel metal2 s 213090 0 213146 800 6 wb_dat_o[23]
port 88 nsew signal output
rlabel metal2 s 221370 0 221426 800 6 wb_dat_o[24]
port 89 nsew signal output
rlabel metal2 s 229558 0 229614 800 6 wb_dat_o[25]
port 90 nsew signal output
rlabel metal2 s 237838 0 237894 800 6 wb_dat_o[26]
port 91 nsew signal output
rlabel metal2 s 246118 0 246174 800 6 wb_dat_o[27]
port 92 nsew signal output
rlabel metal2 s 254398 0 254454 800 6 wb_dat_o[28]
port 93 nsew signal output
rlabel metal2 s 262586 0 262642 800 6 wb_dat_o[29]
port 94 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 wb_dat_o[2]
port 95 nsew signal output
rlabel metal2 s 270866 0 270922 800 6 wb_dat_o[30]
port 96 nsew signal output
rlabel metal2 s 279146 0 279202 800 6 wb_dat_o[31]
port 97 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 wb_dat_o[3]
port 98 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 wb_dat_o[4]
port 99 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 wb_dat_o[5]
port 100 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 wb_dat_o[6]
port 101 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 wb_dat_o[7]
port 102 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 wb_dat_o[8]
port 103 nsew signal output
rlabel metal2 s 97538 0 97594 800 6 wb_dat_o[9]
port 104 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 wb_rst_i
port 105 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wb_stb_i
port 106 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wb_we_i
port 107 nsew signal input
rlabel metal3 s 282526 6672 283326 6792 6 x[0]
port 108 nsew signal input
rlabel metal3 s 282526 141040 283326 141160 6 x[10]
port 109 nsew signal input
rlabel metal3 s 282526 154504 283326 154624 6 x[11]
port 110 nsew signal input
rlabel metal3 s 282526 167968 283326 168088 6 x[12]
port 111 nsew signal input
rlabel metal3 s 282526 181432 283326 181552 6 x[13]
port 112 nsew signal input
rlabel metal3 s 282526 194896 283326 195016 6 x[14]
port 113 nsew signal input
rlabel metal3 s 282526 208360 283326 208480 6 x[15]
port 114 nsew signal input
rlabel metal3 s 282526 20000 283326 20120 6 x[1]
port 115 nsew signal input
rlabel metal3 s 282526 33464 283326 33584 6 x[2]
port 116 nsew signal input
rlabel metal3 s 282526 46928 283326 47048 6 x[3]
port 117 nsew signal input
rlabel metal3 s 282526 60392 283326 60512 6 x[4]
port 118 nsew signal input
rlabel metal3 s 282526 73856 283326 73976 6 x[5]
port 119 nsew signal input
rlabel metal3 s 282526 87320 283326 87440 6 x[6]
port 120 nsew signal input
rlabel metal3 s 282526 100784 283326 100904 6 x[7]
port 121 nsew signal input
rlabel metal3 s 282526 114248 283326 114368 6 x[8]
port 122 nsew signal input
rlabel metal3 s 282526 127576 283326 127696 6 x[9]
port 123 nsew signal input
rlabel metal2 s 39302 214390 39358 215190 6 y[0]
port 124 nsew signal output
rlabel metal2 s 196714 214390 196770 215190 6 y[10]
port 125 nsew signal output
rlabel metal2 s 212446 214390 212502 215190 6 y[11]
port 126 nsew signal output
rlabel metal2 s 228178 214390 228234 215190 6 y[12]
port 127 nsew signal output
rlabel metal2 s 243910 214390 243966 215190 6 y[13]
port 128 nsew signal output
rlabel metal2 s 259642 214390 259698 215190 6 y[14]
port 129 nsew signal output
rlabel metal2 s 275374 214390 275430 215190 6 y[15]
port 130 nsew signal output
rlabel metal2 s 55034 214390 55090 215190 6 y[1]
port 131 nsew signal output
rlabel metal2 s 70766 214390 70822 215190 6 y[2]
port 132 nsew signal output
rlabel metal2 s 86498 214390 86554 215190 6 y[3]
port 133 nsew signal output
rlabel metal2 s 102230 214390 102286 215190 6 y[4]
port 134 nsew signal output
rlabel metal2 s 117962 214390 118018 215190 6 y[5]
port 135 nsew signal output
rlabel metal2 s 133694 214390 133750 215190 6 y[6]
port 136 nsew signal output
rlabel metal2 s 149518 214390 149574 215190 6 y[7]
port 137 nsew signal output
rlabel metal2 s 165250 214390 165306 215190 6 y[8]
port 138 nsew signal output
rlabel metal2 s 180982 214390 181038 215190 6 y[9]
port 139 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 283326 215190
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 75887290
string GDS_FILE /home/openpdk/caravel/fct-iot-node-project/openlane/bqmain/runs/bqmain/results/finishing/bqmain.magic.gds
string GDS_START 1849152
<< end >>

