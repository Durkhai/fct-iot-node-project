VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO biquad
  CLASS BLOCK ;
  FOREIGN biquad ;
  ORIGIN 0.000 0.000 ;
  SIZE 374.375 BY 385.095 ;
  PIN a11[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END a11[0]
  PIN a11[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 25.200 374.375 25.800 ;
    END
  END a11[1]
  PIN a11[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 60.560 374.375 61.160 ;
    END
  END a11[2]
  PIN a11[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 381.095 112.610 385.095 ;
    END
  END a11[3]
  PIN a11[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END a11[4]
  PIN a11[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 182.960 374.375 183.560 ;
    END
  END a11[5]
  PIN a11[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END a11[6]
  PIN a11[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END a11[7]
  PIN a11[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END a11[8]
  PIN a11[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END a11[9]
  PIN a12[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END a12[0]
  PIN a12[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 381.095 37.630 385.095 ;
    END
  END a12[1]
  PIN a12[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 77.560 374.375 78.160 ;
    END
  END a12[2]
  PIN a12[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 381.095 137.450 385.095 ;
    END
  END a12[3]
  PIN a12[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END a12[4]
  PIN a12[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 200.640 374.375 201.240 ;
    END
  END a12[5]
  PIN a12[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 235.320 374.375 235.920 ;
    END
  END a12[6]
  PIN a12[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END a12[7]
  PIN a12[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 381.095 286.950 385.095 ;
    END
  END a12[8]
  PIN a12[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END a12[9]
  PIN b10[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END b10[0]
  PIN b10[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 381.095 62.470 385.095 ;
    END
  END b10[1]
  PIN b10[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END b10[2]
  PIN b10[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END b10[3]
  PIN b10[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END b10[4]
  PIN b10[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END b10[5]
  PIN b10[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 381.095 237.270 385.095 ;
    END
  END b10[6]
  PIN b10[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 287.680 374.375 288.280 ;
    END
  END b10[7]
  PIN b10[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END b10[8]
  PIN b10[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 357.720 374.375 358.320 ;
    END
  END b10[9]
  PIN b11[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END b11[0]
  PIN b11[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END b11[1]
  PIN b11[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 95.240 374.375 95.840 ;
    END
  END b11[2]
  PIN b11[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END b11[3]
  PIN b11[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 147.600 374.375 148.200 ;
    END
  END b11[4]
  PIN b11[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 381.095 187.130 385.095 ;
    END
  END b11[5]
  PIN b11[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END b11[6]
  PIN b11[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END b11[7]
  PIN b11[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 381.095 312.250 385.095 ;
    END
  END b11[8]
  PIN b11[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 375.400 374.375 376.000 ;
    END
  END b11[9]
  PIN b12[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END b12[0]
  PIN b12[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END b12[1]
  PIN b12[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END b12[2]
  PIN b12[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END b12[3]
  PIN b12[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 165.280 374.375 165.880 ;
    END
  END b12[4]
  PIN b12[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 381.095 212.430 385.095 ;
    END
  END b12[5]
  PIN b12[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 4.000 ;
    END
  END b12[6]
  PIN b12[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END b12[7]
  PIN b12[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END b12[8]
  PIN b12[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 381.095 337.090 385.095 ;
    END
  END b12[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 381.095 12.790 385.095 ;
    END
  END clk
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END enable
  PIN nreset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END nreset
  PIN valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END valid
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 372.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 372.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 372.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 372.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 372.880 ;
    END
  END vssd1
  PIN x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 381.095 87.310 385.095 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 112.920 374.375 113.520 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 217.640 374.375 218.240 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 253.000 374.375 253.600 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 305.360 374.375 305.960 ;
    END
  END x[7]
  PIN x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 323.040 374.375 323.640 ;
    END
  END x[8]
  PIN x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 381.095 361.930 385.095 ;
    END
  END x[9]
  PIN yout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 8.200 374.375 8.800 ;
    END
  END yout[0]
  PIN yout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 42.880 374.375 43.480 ;
    END
  END yout[1]
  PIN yout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 130.600 374.375 131.200 ;
    END
  END yout[2]
  PIN yout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END yout[3]
  PIN yout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 381.095 162.290 385.095 ;
    END
  END yout[4]
  PIN yout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END yout[5]
  PIN yout[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 270.000 374.375 270.600 ;
    END
  END yout[6]
  PIN yout[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 381.095 262.110 385.095 ;
    END
  END yout[7]
  PIN yout[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370.375 340.040 374.375 340.640 ;
    END
  END yout[8]
  PIN yout[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 0.000 363.310 4.000 ;
    END
  END yout[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 368.460 372.725 ;
      LAYER met1 ;
        RECT 5.520 9.280 368.460 372.880 ;
      LAYER met2 ;
        RECT 6.990 380.815 12.230 381.890 ;
        RECT 13.070 380.815 37.070 381.890 ;
        RECT 37.910 380.815 61.910 381.890 ;
        RECT 62.750 380.815 86.750 381.890 ;
        RECT 87.590 380.815 112.050 381.890 ;
        RECT 112.890 380.815 136.890 381.890 ;
        RECT 137.730 380.815 161.730 381.890 ;
        RECT 162.570 380.815 186.570 381.890 ;
        RECT 187.410 380.815 211.870 381.890 ;
        RECT 212.710 380.815 236.710 381.890 ;
        RECT 237.550 380.815 261.550 381.890 ;
        RECT 262.390 380.815 286.390 381.890 ;
        RECT 287.230 380.815 311.690 381.890 ;
        RECT 312.530 380.815 336.530 381.890 ;
        RECT 337.370 380.815 361.370 381.890 ;
        RECT 362.210 380.815 365.610 381.890 ;
        RECT 6.990 4.280 365.610 380.815 ;
        RECT 6.990 3.670 10.390 4.280 ;
        RECT 11.230 3.670 32.010 4.280 ;
        RECT 32.850 3.670 54.090 4.280 ;
        RECT 54.930 3.670 76.170 4.280 ;
        RECT 77.010 3.670 98.250 4.280 ;
        RECT 99.090 3.670 120.330 4.280 ;
        RECT 121.170 3.670 142.410 4.280 ;
        RECT 143.250 3.670 164.490 4.280 ;
        RECT 165.330 3.670 186.570 4.280 ;
        RECT 187.410 3.670 208.190 4.280 ;
        RECT 209.030 3.670 230.270 4.280 ;
        RECT 231.110 3.670 252.350 4.280 ;
        RECT 253.190 3.670 274.430 4.280 ;
        RECT 275.270 3.670 296.510 4.280 ;
        RECT 297.350 3.670 318.590 4.280 ;
        RECT 319.430 3.670 340.670 4.280 ;
        RECT 341.510 3.670 362.750 4.280 ;
        RECT 363.590 3.670 365.610 4.280 ;
      LAYER met3 ;
        RECT 4.000 375.720 369.975 375.865 ;
        RECT 4.400 375.000 369.975 375.720 ;
        RECT 4.400 374.320 370.375 375.000 ;
        RECT 4.000 358.720 370.375 374.320 ;
        RECT 4.000 357.320 369.975 358.720 ;
        RECT 4.000 356.680 370.375 357.320 ;
        RECT 4.400 355.280 370.375 356.680 ;
        RECT 4.000 341.040 370.375 355.280 ;
        RECT 4.000 339.640 369.975 341.040 ;
        RECT 4.000 337.640 370.375 339.640 ;
        RECT 4.400 336.240 370.375 337.640 ;
        RECT 4.000 324.040 370.375 336.240 ;
        RECT 4.000 322.640 369.975 324.040 ;
        RECT 4.000 317.920 370.375 322.640 ;
        RECT 4.400 316.520 370.375 317.920 ;
        RECT 4.000 306.360 370.375 316.520 ;
        RECT 4.000 304.960 369.975 306.360 ;
        RECT 4.000 298.880 370.375 304.960 ;
        RECT 4.400 297.480 370.375 298.880 ;
        RECT 4.000 288.680 370.375 297.480 ;
        RECT 4.000 287.280 369.975 288.680 ;
        RECT 4.000 279.840 370.375 287.280 ;
        RECT 4.400 278.440 370.375 279.840 ;
        RECT 4.000 271.000 370.375 278.440 ;
        RECT 4.000 269.600 369.975 271.000 ;
        RECT 4.000 260.120 370.375 269.600 ;
        RECT 4.400 258.720 370.375 260.120 ;
        RECT 4.000 254.000 370.375 258.720 ;
        RECT 4.000 252.600 369.975 254.000 ;
        RECT 4.000 241.080 370.375 252.600 ;
        RECT 4.400 239.680 370.375 241.080 ;
        RECT 4.000 236.320 370.375 239.680 ;
        RECT 4.000 234.920 369.975 236.320 ;
        RECT 4.000 222.040 370.375 234.920 ;
        RECT 4.400 220.640 370.375 222.040 ;
        RECT 4.000 218.640 370.375 220.640 ;
        RECT 4.000 217.240 369.975 218.640 ;
        RECT 4.000 203.000 370.375 217.240 ;
        RECT 4.400 201.640 370.375 203.000 ;
        RECT 4.400 201.600 369.975 201.640 ;
        RECT 4.000 200.240 369.975 201.600 ;
        RECT 4.000 183.960 370.375 200.240 ;
        RECT 4.000 183.280 369.975 183.960 ;
        RECT 4.400 182.560 369.975 183.280 ;
        RECT 4.400 181.880 370.375 182.560 ;
        RECT 4.000 166.280 370.375 181.880 ;
        RECT 4.000 164.880 369.975 166.280 ;
        RECT 4.000 164.240 370.375 164.880 ;
        RECT 4.400 162.840 370.375 164.240 ;
        RECT 4.000 148.600 370.375 162.840 ;
        RECT 4.000 147.200 369.975 148.600 ;
        RECT 4.000 145.200 370.375 147.200 ;
        RECT 4.400 143.800 370.375 145.200 ;
        RECT 4.000 131.600 370.375 143.800 ;
        RECT 4.000 130.200 369.975 131.600 ;
        RECT 4.000 125.480 370.375 130.200 ;
        RECT 4.400 124.080 370.375 125.480 ;
        RECT 4.000 113.920 370.375 124.080 ;
        RECT 4.000 112.520 369.975 113.920 ;
        RECT 4.000 106.440 370.375 112.520 ;
        RECT 4.400 105.040 370.375 106.440 ;
        RECT 4.000 96.240 370.375 105.040 ;
        RECT 4.000 94.840 369.975 96.240 ;
        RECT 4.000 87.400 370.375 94.840 ;
        RECT 4.400 86.000 370.375 87.400 ;
        RECT 4.000 78.560 370.375 86.000 ;
        RECT 4.000 77.160 369.975 78.560 ;
        RECT 4.000 67.680 370.375 77.160 ;
        RECT 4.400 66.280 370.375 67.680 ;
        RECT 4.000 61.560 370.375 66.280 ;
        RECT 4.000 60.160 369.975 61.560 ;
        RECT 4.000 48.640 370.375 60.160 ;
        RECT 4.400 47.240 370.375 48.640 ;
        RECT 4.000 43.880 370.375 47.240 ;
        RECT 4.000 42.480 369.975 43.880 ;
        RECT 4.000 29.600 370.375 42.480 ;
        RECT 4.400 28.200 370.375 29.600 ;
        RECT 4.000 26.200 370.375 28.200 ;
        RECT 4.000 24.800 369.975 26.200 ;
        RECT 4.000 10.560 370.375 24.800 ;
        RECT 4.400 9.200 370.375 10.560 ;
        RECT 4.400 9.160 369.975 9.200 ;
        RECT 4.000 8.335 369.975 9.160 ;
      LAYER met4 ;
        RECT 47.215 11.735 97.440 371.105 ;
        RECT 99.840 11.735 174.240 371.105 ;
        RECT 176.640 11.735 251.040 371.105 ;
        RECT 253.440 11.735 327.840 371.105 ;
        RECT 330.240 11.735 364.025 371.105 ;
  END
END biquad
END LIBRARY

