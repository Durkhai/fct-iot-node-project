VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO coefio
  CLASS BLOCK ;
  FOREIGN coefio ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN a11[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 596.000 22.450 600.000 ;
    END
  END a11[0]
  PIN a11[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 210.160 900.000 210.760 ;
    END
  END a11[10]
  PIN a11[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 596.000 317.310 600.000 ;
    END
  END a11[11]
  PIN a11[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END a11[12]
  PIN a11[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 257.080 900.000 257.680 ;
    END
  END a11[13]
  PIN a11[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END a11[14]
  PIN a11[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 304.000 900.000 304.600 ;
    END
  END a11[15]
  PIN a11[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 312.840 900.000 313.440 ;
    END
  END a11[16]
  PIN a11[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 0.000 533.510 4.000 ;
    END
  END a11[17]
  PIN a11[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 369.280 900.000 369.880 ;
    END
  END a11[18]
  PIN a11[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END a11[19]
  PIN a11[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END a11[1]
  PIN a11[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END a11[20]
  PIN a11[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 596.000 523.850 600.000 ;
    END
  END a11[21]
  PIN a11[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END a11[22]
  PIN a11[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 481.480 900.000 482.080 ;
    END
  END a11[23]
  PIN a11[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END a11[24]
  PIN a11[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END a11[25]
  PIN a11[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END a11[26]
  PIN a11[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END a11[27]
  PIN a11[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 565.800 900.000 566.400 ;
    END
  END a11[28]
  PIN a11[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 596.000 775.010 600.000 ;
    END
  END a11[29]
  PIN a11[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END a11[2]
  PIN a11[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 0.000 838.030 4.000 ;
    END
  END a11[30]
  PIN a11[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END a11[31]
  PIN a11[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END a11[3]
  PIN a11[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END a11[4]
  PIN a11[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 134.680 900.000 135.280 ;
    END
  END a11[5]
  PIN a11[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END a11[6]
  PIN a11[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END a11[7]
  PIN a11[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END a11[8]
  PIN a11[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END a11[9]
  PIN a12[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END a12[0]
  PIN a12[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END a12[10]
  PIN a12[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 596.000 332.030 600.000 ;
    END
  END a12[11]
  PIN a12[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 238.040 900.000 238.640 ;
    END
  END a12[12]
  PIN a12[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END a12[13]
  PIN a12[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END a12[14]
  PIN a12[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END a12[15]
  PIN a12[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 322.360 900.000 322.960 ;
    END
  END a12[16]
  PIN a12[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 341.400 900.000 342.000 ;
    END
  END a12[17]
  PIN a12[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END a12[18]
  PIN a12[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 596.000 509.130 600.000 ;
    END
  END a12[19]
  PIN a12[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 22.480 900.000 23.080 ;
    END
  END a12[1]
  PIN a12[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 0.000 643.910 4.000 ;
    END
  END a12[20]
  PIN a12[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 416.200 900.000 416.800 ;
    END
  END a12[21]
  PIN a12[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END a12[22]
  PIN a12[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.000 4.000 508.600 ;
    END
  END a12[23]
  PIN a12[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 491.000 900.000 491.600 ;
    END
  END a12[24]
  PIN a12[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 518.880 900.000 519.480 ;
    END
  END a12[25]
  PIN a12[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 537.920 900.000 538.520 ;
    END
  END a12[26]
  PIN a12[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.350 0.000 796.630 4.000 ;
    END
  END a12[27]
  PIN a12[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.670 596.000 700.950 600.000 ;
    END
  END a12[28]
  PIN a12[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END a12[29]
  PIN a12[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 50.360 900.000 50.960 ;
    END
  END a12[2]
  PIN a12[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END a12[30]
  PIN a12[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 596.000 863.330 600.000 ;
    END
  END a12[31]
  PIN a12[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 78.920 900.000 79.520 ;
    END
  END a12[3]
  PIN a12[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 596.000 169.650 600.000 ;
    END
  END a12[4]
  PIN a12[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END a12[5]
  PIN a12[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 144.200 900.000 144.800 ;
    END
  END a12[6]
  PIN a12[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END a12[7]
  PIN a12[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END a12[8]
  PIN a12[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 181.600 900.000 182.200 ;
    END
  END a12[9]
  PIN ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 596.000 7.730 600.000 ;
    END
  END ack_o
  PIN adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 596.000 37.170 600.000 ;
    END
  END adr_i[0]
  PIN adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 32.000 900.000 32.600 ;
    END
  END adr_i[1]
  PIN adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 59.880 900.000 60.480 ;
    END
  END adr_i[2]
  PIN adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END adr_i[3]
  PIN b10[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END b10[0]
  PIN b10[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END b10[10]
  PIN b10[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 596.000 346.750 600.000 ;
    END
  END b10[11]
  PIN b10[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END b10[12]
  PIN b10[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 596.000 376.650 600.000 ;
    END
  END b10[13]
  PIN b10[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 596.000 391.370 600.000 ;
    END
  END b10[14]
  PIN b10[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END b10[15]
  PIN b10[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 596.000 435.530 600.000 ;
    END
  END b10[16]
  PIN b10[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 596.000 479.690 600.000 ;
    END
  END b10[17]
  PIN b10[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 0.000 588.710 4.000 ;
    END
  END b10[18]
  PIN b10[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 0.000 616.310 4.000 ;
    END
  END b10[19]
  PIN b10[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 41.520 900.000 42.120 ;
    END
  END b10[1]
  PIN b10[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END b10[20]
  PIN b10[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 425.720 900.000 426.320 ;
    END
  END b10[21]
  PIN b10[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END b10[22]
  PIN b10[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END b10[23]
  PIN b10[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END b10[24]
  PIN b10[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 596.000 612.630 600.000 ;
    END
  END b10[25]
  PIN b10[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 0.000 754.770 4.000 ;
    END
  END b10[26]
  PIN b10[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 0.000 810.430 4.000 ;
    END
  END b10[27]
  PIN b10[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 596.000 715.670 600.000 ;
    END
  END b10[28]
  PIN b10[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 584.840 900.000 585.440 ;
    END
  END b10[29]
  PIN b10[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END b10[2]
  PIN b10[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.550 0.000 851.830 4.000 ;
    END
  END b10[30]
  PIN b10[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END b10[31]
  PIN b10[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 88.440 900.000 89.040 ;
    END
  END b10[3]
  PIN b10[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 116.320 900.000 116.920 ;
    END
  END b10[4]
  PIN b10[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END b10[5]
  PIN b10[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END b10[6]
  PIN b10[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END b10[7]
  PIN b10[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END b10[8]
  PIN b10[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END b10[9]
  PIN b11[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END b11[0]
  PIN b11[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END b11[10]
  PIN b11[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END b11[11]
  PIN b11[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END b11[12]
  PIN b11[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END b11[13]
  PIN b11[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 284.960 900.000 285.560 ;
    END
  END b11[14]
  PIN b11[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 596.000 406.090 600.000 ;
    END
  END b11[15]
  PIN b11[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END b11[16]
  PIN b11[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 350.240 900.000 350.840 ;
    END
  END b11[17]
  PIN b11[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.280 4.000 437.880 ;
    END
  END b11[18]
  PIN b11[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END b11[19]
  PIN b11[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END b11[1]
  PIN b11[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END b11[20]
  PIN b11[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 434.560 900.000 435.160 ;
    END
  END b11[21]
  PIN b11[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 596.000 538.570 600.000 ;
    END
  END b11[22]
  PIN b11[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.160 4.000 516.760 ;
    END
  END b11[23]
  PIN b11[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 500.520 900.000 501.120 ;
    END
  END b11[24]
  PIN b11[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.070 596.000 627.350 600.000 ;
    END
  END b11[25]
  PIN b11[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 547.440 900.000 548.040 ;
    END
  END b11[26]
  PIN b11[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 596.000 671.510 600.000 ;
    END
  END b11[27]
  PIN b11[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 596.000 730.850 600.000 ;
    END
  END b11[28]
  PIN b11[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 596.000 789.730 600.000 ;
    END
  END b11[29]
  PIN b11[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END b11[2]
  PIN b11[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END b11[30]
  PIN b11[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 594.360 900.000 594.960 ;
    END
  END b11[31]
  PIN b11[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 596.000 125.490 600.000 ;
    END
  END b11[3]
  PIN b11[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END b11[4]
  PIN b11[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 596.000 199.550 600.000 ;
    END
  END b11[5]
  PIN b11[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END b11[6]
  PIN b11[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 153.720 900.000 154.320 ;
    END
  END b11[7]
  PIN b11[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END b11[8]
  PIN b11[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 191.120 900.000 191.720 ;
    END
  END b11[9]
  PIN b12[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END b12[0]
  PIN b12[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 4.000 ;
    END
  END b12[10]
  PIN b12[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END b12[11]
  PIN b12[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 596.000 361.470 600.000 ;
    END
  END b12[12]
  PIN b12[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 265.920 900.000 266.520 ;
    END
  END b12[13]
  PIN b12[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END b12[14]
  PIN b12[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 596.000 420.810 600.000 ;
    END
  END b12[15]
  PIN b12[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 596.000 450.250 600.000 ;
    END
  END b12[16]
  PIN b12[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 0.000 547.310 4.000 ;
    END
  END b12[17]
  PIN b12[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 596.000 494.410 600.000 ;
    END
  END b12[18]
  PIN b12[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 388.320 900.000 388.920 ;
    END
  END b12[19]
  PIN b12[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END b12[1]
  PIN b12[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 4.000 ;
    END
  END b12[20]
  PIN b12[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 444.080 900.000 444.680 ;
    END
  END b12[21]
  PIN b12[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 596.000 553.750 600.000 ;
    END
  END b12[22]
  PIN b12[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 596.000 568.470 600.000 ;
    END
  END b12[23]
  PIN b12[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 0.000 727.170 4.000 ;
    END
  END b12[24]
  PIN b12[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 596.000 642.070 600.000 ;
    END
  END b12[25]
  PIN b12[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 556.960 900.000 557.560 ;
    END
  END b12[26]
  PIN b12[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 596.000 686.230 600.000 ;
    END
  END b12[27]
  PIN b12[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 596.000 745.570 600.000 ;
    END
  END b12[28]
  PIN b12[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 596.000 804.450 600.000 ;
    END
  END b12[29]
  PIN b12[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END b12[2]
  PIN b12[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.880 4.000 587.480 ;
    END
  END b12[30]
  PIN b12[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.950 0.000 893.230 4.000 ;
    END
  END b12[31]
  PIN b12[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 596.000 140.210 600.000 ;
    END
  END b12[3]
  PIN b12[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END b12[4]
  PIN b12[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END b12[5]
  PIN b12[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END b12[6]
  PIN b12[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 596.000 273.150 600.000 ;
    END
  END b12[7]
  PIN b12[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END b12[8]
  PIN b12[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 596.000 302.590 600.000 ;
    END
  END b12[9]
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END clk_i
  PIN cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END cyc_i
  PIN dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END dat_i[0]
  PIN dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END dat_i[10]
  PIN dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 219.000 900.000 219.600 ;
    END
  END dat_i[11]
  PIN dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END dat_i[12]
  PIN dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END dat_i[13]
  PIN dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END dat_i[14]
  PIN dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END dat_i[15]
  PIN dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 596.000 464.970 600.000 ;
    END
  END dat_i[16]
  PIN dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 359.760 900.000 360.360 ;
    END
  END dat_i[17]
  PIN dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 378.800 900.000 379.400 ;
    END
  END dat_i[18]
  PIN dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 0.000 630.110 4.000 ;
    END
  END dat_i[19]
  PIN dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 596.000 81.330 600.000 ;
    END
  END dat_i[1]
  PIN dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 406.680 900.000 407.280 ;
    END
  END dat_i[20]
  PIN dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 453.600 900.000 454.200 ;
    END
  END dat_i[21]
  PIN dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 463.120 900.000 463.720 ;
    END
  END dat_i[22]
  PIN dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 596.000 583.190 600.000 ;
    END
  END dat_i[23]
  PIN dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 596.000 597.910 600.000 ;
    END
  END dat_i[24]
  PIN dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 528.400 900.000 529.000 ;
    END
  END dat_i[25]
  PIN dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 596.000 656.790 600.000 ;
    END
  END dat_i[26]
  PIN dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 0.000 824.230 4.000 ;
    END
  END dat_i[27]
  PIN dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 596.000 760.290 600.000 ;
    END
  END dat_i[28]
  PIN dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 596.000 819.170 600.000 ;
    END
  END dat_i[29]
  PIN dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 69.400 900.000 70.000 ;
    END
  END dat_i[2]
  PIN dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 596.000 848.610 600.000 ;
    END
  END dat_i[30]
  PIN dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 596.000 878.050 600.000 ;
    END
  END dat_i[31]
  PIN dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 596.000 154.930 600.000 ;
    END
  END dat_i[3]
  PIN dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 4.000 145.480 ;
    END
  END dat_i[4]
  PIN dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END dat_i[5]
  PIN dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END dat_i[6]
  PIN dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END dat_i[7]
  PIN dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 163.240 900.000 163.840 ;
    END
  END dat_i[8]
  PIN dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END dat_i[9]
  PIN dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 596.000 51.890 600.000 ;
    END
  END dat_o[0]
  PIN dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END dat_o[10]
  PIN dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 228.520 900.000 229.120 ;
    END
  END dat_o[11]
  PIN dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END dat_o[12]
  PIN dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END dat_o[13]
  PIN dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 0.000 477.850 4.000 ;
    END
  END dat_o[14]
  PIN dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 0.000 519.250 4.000 ;
    END
  END dat_o[15]
  PIN dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 331.880 900.000 332.480 ;
    END
  END dat_o[16]
  PIN dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 4.000 ;
    END
  END dat_o[17]
  PIN dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END dat_o[18]
  PIN dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 397.160 900.000 397.760 ;
    END
  END dat_o[19]
  PIN dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END dat_o[1]
  PIN dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END dat_o[20]
  PIN dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END dat_o[21]
  PIN dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 472.640 900.000 473.240 ;
    END
  END dat_o[22]
  PIN dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 0.000 713.370 4.000 ;
    END
  END dat_o[23]
  PIN dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 510.040 900.000 510.640 ;
    END
  END dat_o[24]
  PIN dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END dat_o[25]
  PIN dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 4.000 ;
    END
  END dat_o[26]
  PIN dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 555.600 4.000 556.200 ;
    END
  END dat_o[27]
  PIN dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 575.320 900.000 575.920 ;
    END
  END dat_o[28]
  PIN dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.610 596.000 833.890 600.000 ;
    END
  END dat_o[29]
  PIN dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 596.000 110.770 600.000 ;
    END
  END dat_o[2]
  PIN dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.350 0.000 865.630 4.000 ;
    END
  END dat_o[30]
  PIN dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 596.000 892.770 600.000 ;
    END
  END dat_o[31]
  PIN dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 97.280 900.000 97.880 ;
    END
  END dat_o[3]
  PIN dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 596.000 184.370 600.000 ;
    END
  END dat_o[4]
  PIN dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 596.000 214.270 600.000 ;
    END
  END dat_o[5]
  PIN dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 596.000 258.430 600.000 ;
    END
  END dat_o[6]
  PIN dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END dat_o[7]
  PIN dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 172.760 900.000 173.360 ;
    END
  END dat_o[8]
  PIN dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END dat_o[9]
  PIN rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 4.120 900.000 4.720 ;
    END
  END rst_i
  PIN stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 12.960 900.000 13.560 ;
    END
  END stb_i
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END we_i
  PIN x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 596.000 66.610 600.000 ;
    END
  END x[0]
  PIN x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END x[10]
  PIN x[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.960 4.000 319.560 ;
    END
  END x[11]
  PIN x[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 247.560 900.000 248.160 ;
    END
  END x[12]
  PIN x[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END x[13]
  PIN x[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 294.480 900.000 295.080 ;
    END
  END x[14]
  PIN x[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END x[15]
  PIN x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 125.840 900.000 126.440 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 596.000 228.990 600.000 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 596.000 287.870 600.000 ;
    END
  END x[7]
  PIN x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END x[8]
  PIN x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END x[9]
  PIN y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END y[0]
  PIN y[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END y[10]
  PIN y[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END y[11]
  PIN y[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END y[12]
  PIN y[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 275.440 900.000 276.040 ;
    END
  END y[13]
  PIN y[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END y[14]
  PIN y[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END y[15]
  PIN y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 596.000 96.050 600.000 ;
    END
  END y[1]
  PIN y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END y[2]
  PIN y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 106.800 900.000 107.400 ;
    END
  END y[3]
  PIN y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END y[4]
  PIN y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 596.000 243.710 600.000 ;
    END
  END y[5]
  PIN y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END y[6]
  PIN y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END y[7]
  PIN y[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END y[8]
  PIN y[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 200.640 900.000 201.240 ;
    END
  END y[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 9.900 894.240 587.760 ;
      LAYER met2 ;
        RECT 6.990 595.720 7.170 596.770 ;
        RECT 8.010 595.720 21.890 596.770 ;
        RECT 22.730 595.720 36.610 596.770 ;
        RECT 37.450 595.720 51.330 596.770 ;
        RECT 52.170 595.720 66.050 596.770 ;
        RECT 66.890 595.720 80.770 596.770 ;
        RECT 81.610 595.720 95.490 596.770 ;
        RECT 96.330 595.720 110.210 596.770 ;
        RECT 111.050 595.720 124.930 596.770 ;
        RECT 125.770 595.720 139.650 596.770 ;
        RECT 140.490 595.720 154.370 596.770 ;
        RECT 155.210 595.720 169.090 596.770 ;
        RECT 169.930 595.720 183.810 596.770 ;
        RECT 184.650 595.720 198.990 596.770 ;
        RECT 199.830 595.720 213.710 596.770 ;
        RECT 214.550 595.720 228.430 596.770 ;
        RECT 229.270 595.720 243.150 596.770 ;
        RECT 243.990 595.720 257.870 596.770 ;
        RECT 258.710 595.720 272.590 596.770 ;
        RECT 273.430 595.720 287.310 596.770 ;
        RECT 288.150 595.720 302.030 596.770 ;
        RECT 302.870 595.720 316.750 596.770 ;
        RECT 317.590 595.720 331.470 596.770 ;
        RECT 332.310 595.720 346.190 596.770 ;
        RECT 347.030 595.720 360.910 596.770 ;
        RECT 361.750 595.720 376.090 596.770 ;
        RECT 376.930 595.720 390.810 596.770 ;
        RECT 391.650 595.720 405.530 596.770 ;
        RECT 406.370 595.720 420.250 596.770 ;
        RECT 421.090 595.720 434.970 596.770 ;
        RECT 435.810 595.720 449.690 596.770 ;
        RECT 450.530 595.720 464.410 596.770 ;
        RECT 465.250 595.720 479.130 596.770 ;
        RECT 479.970 595.720 493.850 596.770 ;
        RECT 494.690 595.720 508.570 596.770 ;
        RECT 509.410 595.720 523.290 596.770 ;
        RECT 524.130 595.720 538.010 596.770 ;
        RECT 538.850 595.720 553.190 596.770 ;
        RECT 554.030 595.720 567.910 596.770 ;
        RECT 568.750 595.720 582.630 596.770 ;
        RECT 583.470 595.720 597.350 596.770 ;
        RECT 598.190 595.720 612.070 596.770 ;
        RECT 612.910 595.720 626.790 596.770 ;
        RECT 627.630 595.720 641.510 596.770 ;
        RECT 642.350 595.720 656.230 596.770 ;
        RECT 657.070 595.720 670.950 596.770 ;
        RECT 671.790 595.720 685.670 596.770 ;
        RECT 686.510 595.720 700.390 596.770 ;
        RECT 701.230 595.720 715.110 596.770 ;
        RECT 715.950 595.720 730.290 596.770 ;
        RECT 731.130 595.720 745.010 596.770 ;
        RECT 745.850 595.720 759.730 596.770 ;
        RECT 760.570 595.720 774.450 596.770 ;
        RECT 775.290 595.720 789.170 596.770 ;
        RECT 790.010 595.720 803.890 596.770 ;
        RECT 804.730 595.720 818.610 596.770 ;
        RECT 819.450 595.720 833.330 596.770 ;
        RECT 834.170 595.720 848.050 596.770 ;
        RECT 848.890 595.720 862.770 596.770 ;
        RECT 863.610 595.720 877.490 596.770 ;
        RECT 878.330 595.720 892.210 596.770 ;
        RECT 893.050 595.720 893.220 596.770 ;
        RECT 6.990 4.280 893.220 595.720 ;
        RECT 7.550 3.555 20.510 4.280 ;
        RECT 21.350 3.555 34.310 4.280 ;
        RECT 35.150 3.555 48.110 4.280 ;
        RECT 48.950 3.555 61.910 4.280 ;
        RECT 62.750 3.555 75.710 4.280 ;
        RECT 76.550 3.555 89.510 4.280 ;
        RECT 90.350 3.555 103.310 4.280 ;
        RECT 104.150 3.555 117.110 4.280 ;
        RECT 117.950 3.555 130.910 4.280 ;
        RECT 131.750 3.555 145.170 4.280 ;
        RECT 146.010 3.555 158.970 4.280 ;
        RECT 159.810 3.555 172.770 4.280 ;
        RECT 173.610 3.555 186.570 4.280 ;
        RECT 187.410 3.555 200.370 4.280 ;
        RECT 201.210 3.555 214.170 4.280 ;
        RECT 215.010 3.555 227.970 4.280 ;
        RECT 228.810 3.555 241.770 4.280 ;
        RECT 242.610 3.555 255.570 4.280 ;
        RECT 256.410 3.555 269.830 4.280 ;
        RECT 270.670 3.555 283.630 4.280 ;
        RECT 284.470 3.555 297.430 4.280 ;
        RECT 298.270 3.555 311.230 4.280 ;
        RECT 312.070 3.555 325.030 4.280 ;
        RECT 325.870 3.555 338.830 4.280 ;
        RECT 339.670 3.555 352.630 4.280 ;
        RECT 353.470 3.555 366.430 4.280 ;
        RECT 367.270 3.555 380.230 4.280 ;
        RECT 381.070 3.555 394.490 4.280 ;
        RECT 395.330 3.555 408.290 4.280 ;
        RECT 409.130 3.555 422.090 4.280 ;
        RECT 422.930 3.555 435.890 4.280 ;
        RECT 436.730 3.555 449.690 4.280 ;
        RECT 450.530 3.555 463.490 4.280 ;
        RECT 464.330 3.555 477.290 4.280 ;
        RECT 478.130 3.555 491.090 4.280 ;
        RECT 491.930 3.555 504.890 4.280 ;
        RECT 505.730 3.555 518.690 4.280 ;
        RECT 519.530 3.555 532.950 4.280 ;
        RECT 533.790 3.555 546.750 4.280 ;
        RECT 547.590 3.555 560.550 4.280 ;
        RECT 561.390 3.555 574.350 4.280 ;
        RECT 575.190 3.555 588.150 4.280 ;
        RECT 588.990 3.555 601.950 4.280 ;
        RECT 602.790 3.555 615.750 4.280 ;
        RECT 616.590 3.555 629.550 4.280 ;
        RECT 630.390 3.555 643.350 4.280 ;
        RECT 644.190 3.555 657.610 4.280 ;
        RECT 658.450 3.555 671.410 4.280 ;
        RECT 672.250 3.555 685.210 4.280 ;
        RECT 686.050 3.555 699.010 4.280 ;
        RECT 699.850 3.555 712.810 4.280 ;
        RECT 713.650 3.555 726.610 4.280 ;
        RECT 727.450 3.555 740.410 4.280 ;
        RECT 741.250 3.555 754.210 4.280 ;
        RECT 755.050 3.555 768.010 4.280 ;
        RECT 768.850 3.555 782.270 4.280 ;
        RECT 783.110 3.555 796.070 4.280 ;
        RECT 796.910 3.555 809.870 4.280 ;
        RECT 810.710 3.555 823.670 4.280 ;
        RECT 824.510 3.555 837.470 4.280 ;
        RECT 838.310 3.555 851.270 4.280 ;
        RECT 852.110 3.555 865.070 4.280 ;
        RECT 865.910 3.555 878.870 4.280 ;
        RECT 879.710 3.555 892.670 4.280 ;
      LAYER met3 ;
        RECT 4.400 595.360 896.000 595.505 ;
        RECT 4.400 594.640 895.600 595.360 ;
        RECT 4.000 593.960 895.600 594.640 ;
        RECT 4.000 587.880 896.000 593.960 ;
        RECT 4.400 586.480 896.000 587.880 ;
        RECT 4.000 585.840 896.000 586.480 ;
        RECT 4.000 584.440 895.600 585.840 ;
        RECT 4.000 580.400 896.000 584.440 ;
        RECT 4.400 579.000 896.000 580.400 ;
        RECT 4.000 576.320 896.000 579.000 ;
        RECT 4.000 574.920 895.600 576.320 ;
        RECT 4.000 572.240 896.000 574.920 ;
        RECT 4.400 570.840 896.000 572.240 ;
        RECT 4.000 566.800 896.000 570.840 ;
        RECT 4.000 565.400 895.600 566.800 ;
        RECT 4.000 564.080 896.000 565.400 ;
        RECT 4.400 562.680 896.000 564.080 ;
        RECT 4.000 557.960 896.000 562.680 ;
        RECT 4.000 556.600 895.600 557.960 ;
        RECT 4.400 556.560 895.600 556.600 ;
        RECT 4.400 555.200 896.000 556.560 ;
        RECT 4.000 548.440 896.000 555.200 ;
        RECT 4.400 547.040 895.600 548.440 ;
        RECT 4.000 540.960 896.000 547.040 ;
        RECT 4.400 539.560 896.000 540.960 ;
        RECT 4.000 538.920 896.000 539.560 ;
        RECT 4.000 537.520 895.600 538.920 ;
        RECT 4.000 532.800 896.000 537.520 ;
        RECT 4.400 531.400 896.000 532.800 ;
        RECT 4.000 529.400 896.000 531.400 ;
        RECT 4.000 528.000 895.600 529.400 ;
        RECT 4.000 524.640 896.000 528.000 ;
        RECT 4.400 523.240 896.000 524.640 ;
        RECT 4.000 519.880 896.000 523.240 ;
        RECT 4.000 518.480 895.600 519.880 ;
        RECT 4.000 517.160 896.000 518.480 ;
        RECT 4.400 515.760 896.000 517.160 ;
        RECT 4.000 511.040 896.000 515.760 ;
        RECT 4.000 509.640 895.600 511.040 ;
        RECT 4.000 509.000 896.000 509.640 ;
        RECT 4.400 507.600 896.000 509.000 ;
        RECT 4.000 501.520 896.000 507.600 ;
        RECT 4.400 500.120 895.600 501.520 ;
        RECT 4.000 493.360 896.000 500.120 ;
        RECT 4.400 492.000 896.000 493.360 ;
        RECT 4.400 491.960 895.600 492.000 ;
        RECT 4.000 490.600 895.600 491.960 ;
        RECT 4.000 485.200 896.000 490.600 ;
        RECT 4.400 483.800 896.000 485.200 ;
        RECT 4.000 482.480 896.000 483.800 ;
        RECT 4.000 481.080 895.600 482.480 ;
        RECT 4.000 477.720 896.000 481.080 ;
        RECT 4.400 476.320 896.000 477.720 ;
        RECT 4.000 473.640 896.000 476.320 ;
        RECT 4.000 472.240 895.600 473.640 ;
        RECT 4.000 469.560 896.000 472.240 ;
        RECT 4.400 468.160 896.000 469.560 ;
        RECT 4.000 464.120 896.000 468.160 ;
        RECT 4.000 462.720 895.600 464.120 ;
        RECT 4.000 462.080 896.000 462.720 ;
        RECT 4.400 460.680 896.000 462.080 ;
        RECT 4.000 454.600 896.000 460.680 ;
        RECT 4.000 453.920 895.600 454.600 ;
        RECT 4.400 453.200 895.600 453.920 ;
        RECT 4.400 452.520 896.000 453.200 ;
        RECT 4.000 445.760 896.000 452.520 ;
        RECT 4.400 445.080 896.000 445.760 ;
        RECT 4.400 444.360 895.600 445.080 ;
        RECT 4.000 443.680 895.600 444.360 ;
        RECT 4.000 438.280 896.000 443.680 ;
        RECT 4.400 436.880 896.000 438.280 ;
        RECT 4.000 435.560 896.000 436.880 ;
        RECT 4.000 434.160 895.600 435.560 ;
        RECT 4.000 430.120 896.000 434.160 ;
        RECT 4.400 428.720 896.000 430.120 ;
        RECT 4.000 426.720 896.000 428.720 ;
        RECT 4.000 425.320 895.600 426.720 ;
        RECT 4.000 422.640 896.000 425.320 ;
        RECT 4.400 421.240 896.000 422.640 ;
        RECT 4.000 417.200 896.000 421.240 ;
        RECT 4.000 415.800 895.600 417.200 ;
        RECT 4.000 414.480 896.000 415.800 ;
        RECT 4.400 413.080 896.000 414.480 ;
        RECT 4.000 407.680 896.000 413.080 ;
        RECT 4.000 406.320 895.600 407.680 ;
        RECT 4.400 406.280 895.600 406.320 ;
        RECT 4.400 404.920 896.000 406.280 ;
        RECT 4.000 398.840 896.000 404.920 ;
        RECT 4.400 398.160 896.000 398.840 ;
        RECT 4.400 397.440 895.600 398.160 ;
        RECT 4.000 396.760 895.600 397.440 ;
        RECT 4.000 390.680 896.000 396.760 ;
        RECT 4.400 389.320 896.000 390.680 ;
        RECT 4.400 389.280 895.600 389.320 ;
        RECT 4.000 387.920 895.600 389.280 ;
        RECT 4.000 383.200 896.000 387.920 ;
        RECT 4.400 381.800 896.000 383.200 ;
        RECT 4.000 379.800 896.000 381.800 ;
        RECT 4.000 378.400 895.600 379.800 ;
        RECT 4.000 375.040 896.000 378.400 ;
        RECT 4.400 373.640 896.000 375.040 ;
        RECT 4.000 370.280 896.000 373.640 ;
        RECT 4.000 368.880 895.600 370.280 ;
        RECT 4.000 366.880 896.000 368.880 ;
        RECT 4.400 365.480 896.000 366.880 ;
        RECT 4.000 360.760 896.000 365.480 ;
        RECT 4.000 359.400 895.600 360.760 ;
        RECT 4.400 359.360 895.600 359.400 ;
        RECT 4.400 358.000 896.000 359.360 ;
        RECT 4.000 351.240 896.000 358.000 ;
        RECT 4.400 349.840 895.600 351.240 ;
        RECT 4.000 343.760 896.000 349.840 ;
        RECT 4.400 342.400 896.000 343.760 ;
        RECT 4.400 342.360 895.600 342.400 ;
        RECT 4.000 341.000 895.600 342.360 ;
        RECT 4.000 335.600 896.000 341.000 ;
        RECT 4.400 334.200 896.000 335.600 ;
        RECT 4.000 332.880 896.000 334.200 ;
        RECT 4.000 331.480 895.600 332.880 ;
        RECT 4.000 327.440 896.000 331.480 ;
        RECT 4.400 326.040 896.000 327.440 ;
        RECT 4.000 323.360 896.000 326.040 ;
        RECT 4.000 321.960 895.600 323.360 ;
        RECT 4.000 319.960 896.000 321.960 ;
        RECT 4.400 318.560 896.000 319.960 ;
        RECT 4.000 313.840 896.000 318.560 ;
        RECT 4.000 312.440 895.600 313.840 ;
        RECT 4.000 311.800 896.000 312.440 ;
        RECT 4.400 310.400 896.000 311.800 ;
        RECT 4.000 305.000 896.000 310.400 ;
        RECT 4.000 304.320 895.600 305.000 ;
        RECT 4.400 303.600 895.600 304.320 ;
        RECT 4.400 302.920 896.000 303.600 ;
        RECT 4.000 296.160 896.000 302.920 ;
        RECT 4.400 295.480 896.000 296.160 ;
        RECT 4.400 294.760 895.600 295.480 ;
        RECT 4.000 294.080 895.600 294.760 ;
        RECT 4.000 288.000 896.000 294.080 ;
        RECT 4.400 286.600 896.000 288.000 ;
        RECT 4.000 285.960 896.000 286.600 ;
        RECT 4.000 284.560 895.600 285.960 ;
        RECT 4.000 280.520 896.000 284.560 ;
        RECT 4.400 279.120 896.000 280.520 ;
        RECT 4.000 276.440 896.000 279.120 ;
        RECT 4.000 275.040 895.600 276.440 ;
        RECT 4.000 272.360 896.000 275.040 ;
        RECT 4.400 270.960 896.000 272.360 ;
        RECT 4.000 266.920 896.000 270.960 ;
        RECT 4.000 265.520 895.600 266.920 ;
        RECT 4.000 264.200 896.000 265.520 ;
        RECT 4.400 262.800 896.000 264.200 ;
        RECT 4.000 258.080 896.000 262.800 ;
        RECT 4.000 256.720 895.600 258.080 ;
        RECT 4.400 256.680 895.600 256.720 ;
        RECT 4.400 255.320 896.000 256.680 ;
        RECT 4.000 248.560 896.000 255.320 ;
        RECT 4.400 247.160 895.600 248.560 ;
        RECT 4.000 241.080 896.000 247.160 ;
        RECT 4.400 239.680 896.000 241.080 ;
        RECT 4.000 239.040 896.000 239.680 ;
        RECT 4.000 237.640 895.600 239.040 ;
        RECT 4.000 232.920 896.000 237.640 ;
        RECT 4.400 231.520 896.000 232.920 ;
        RECT 4.000 229.520 896.000 231.520 ;
        RECT 4.000 228.120 895.600 229.520 ;
        RECT 4.000 224.760 896.000 228.120 ;
        RECT 4.400 223.360 896.000 224.760 ;
        RECT 4.000 220.000 896.000 223.360 ;
        RECT 4.000 218.600 895.600 220.000 ;
        RECT 4.000 217.280 896.000 218.600 ;
        RECT 4.400 215.880 896.000 217.280 ;
        RECT 4.000 211.160 896.000 215.880 ;
        RECT 4.000 209.760 895.600 211.160 ;
        RECT 4.000 209.120 896.000 209.760 ;
        RECT 4.400 207.720 896.000 209.120 ;
        RECT 4.000 201.640 896.000 207.720 ;
        RECT 4.400 200.240 895.600 201.640 ;
        RECT 4.000 193.480 896.000 200.240 ;
        RECT 4.400 192.120 896.000 193.480 ;
        RECT 4.400 192.080 895.600 192.120 ;
        RECT 4.000 190.720 895.600 192.080 ;
        RECT 4.000 185.320 896.000 190.720 ;
        RECT 4.400 183.920 896.000 185.320 ;
        RECT 4.000 182.600 896.000 183.920 ;
        RECT 4.000 181.200 895.600 182.600 ;
        RECT 4.000 177.840 896.000 181.200 ;
        RECT 4.400 176.440 896.000 177.840 ;
        RECT 4.000 173.760 896.000 176.440 ;
        RECT 4.000 172.360 895.600 173.760 ;
        RECT 4.000 169.680 896.000 172.360 ;
        RECT 4.400 168.280 896.000 169.680 ;
        RECT 4.000 164.240 896.000 168.280 ;
        RECT 4.000 162.840 895.600 164.240 ;
        RECT 4.000 162.200 896.000 162.840 ;
        RECT 4.400 160.800 896.000 162.200 ;
        RECT 4.000 154.720 896.000 160.800 ;
        RECT 4.000 154.040 895.600 154.720 ;
        RECT 4.400 153.320 895.600 154.040 ;
        RECT 4.400 152.640 896.000 153.320 ;
        RECT 4.000 145.880 896.000 152.640 ;
        RECT 4.400 145.200 896.000 145.880 ;
        RECT 4.400 144.480 895.600 145.200 ;
        RECT 4.000 143.800 895.600 144.480 ;
        RECT 4.000 138.400 896.000 143.800 ;
        RECT 4.400 137.000 896.000 138.400 ;
        RECT 4.000 135.680 896.000 137.000 ;
        RECT 4.000 134.280 895.600 135.680 ;
        RECT 4.000 130.240 896.000 134.280 ;
        RECT 4.400 128.840 896.000 130.240 ;
        RECT 4.000 126.840 896.000 128.840 ;
        RECT 4.000 125.440 895.600 126.840 ;
        RECT 4.000 122.760 896.000 125.440 ;
        RECT 4.400 121.360 896.000 122.760 ;
        RECT 4.000 117.320 896.000 121.360 ;
        RECT 4.000 115.920 895.600 117.320 ;
        RECT 4.000 114.600 896.000 115.920 ;
        RECT 4.400 113.200 896.000 114.600 ;
        RECT 4.000 107.800 896.000 113.200 ;
        RECT 4.000 106.440 895.600 107.800 ;
        RECT 4.400 106.400 895.600 106.440 ;
        RECT 4.400 105.040 896.000 106.400 ;
        RECT 4.000 98.960 896.000 105.040 ;
        RECT 4.400 98.280 896.000 98.960 ;
        RECT 4.400 97.560 895.600 98.280 ;
        RECT 4.000 96.880 895.600 97.560 ;
        RECT 4.000 90.800 896.000 96.880 ;
        RECT 4.400 89.440 896.000 90.800 ;
        RECT 4.400 89.400 895.600 89.440 ;
        RECT 4.000 88.040 895.600 89.400 ;
        RECT 4.000 83.320 896.000 88.040 ;
        RECT 4.400 81.920 896.000 83.320 ;
        RECT 4.000 79.920 896.000 81.920 ;
        RECT 4.000 78.520 895.600 79.920 ;
        RECT 4.000 75.160 896.000 78.520 ;
        RECT 4.400 73.760 896.000 75.160 ;
        RECT 4.000 70.400 896.000 73.760 ;
        RECT 4.000 69.000 895.600 70.400 ;
        RECT 4.000 67.000 896.000 69.000 ;
        RECT 4.400 65.600 896.000 67.000 ;
        RECT 4.000 60.880 896.000 65.600 ;
        RECT 4.000 59.520 895.600 60.880 ;
        RECT 4.400 59.480 895.600 59.520 ;
        RECT 4.400 58.120 896.000 59.480 ;
        RECT 4.000 51.360 896.000 58.120 ;
        RECT 4.400 49.960 895.600 51.360 ;
        RECT 4.000 43.880 896.000 49.960 ;
        RECT 4.400 42.520 896.000 43.880 ;
        RECT 4.400 42.480 895.600 42.520 ;
        RECT 4.000 41.120 895.600 42.480 ;
        RECT 4.000 35.720 896.000 41.120 ;
        RECT 4.400 34.320 896.000 35.720 ;
        RECT 4.000 33.000 896.000 34.320 ;
        RECT 4.000 31.600 895.600 33.000 ;
        RECT 4.000 27.560 896.000 31.600 ;
        RECT 4.400 26.160 896.000 27.560 ;
        RECT 4.000 23.480 896.000 26.160 ;
        RECT 4.000 22.080 895.600 23.480 ;
        RECT 4.000 20.080 896.000 22.080 ;
        RECT 4.400 18.680 896.000 20.080 ;
        RECT 4.000 13.960 896.000 18.680 ;
        RECT 4.000 12.560 895.600 13.960 ;
        RECT 4.000 11.920 896.000 12.560 ;
        RECT 4.400 10.520 896.000 11.920 ;
        RECT 4.000 5.120 896.000 10.520 ;
        RECT 4.000 4.440 895.600 5.120 ;
        RECT 4.400 3.720 895.600 4.440 ;
        RECT 4.400 3.575 896.000 3.720 ;
      LAYER met4 ;
        RECT 285.495 17.175 327.840 569.665 ;
        RECT 330.240 17.175 404.640 569.665 ;
        RECT 407.040 17.175 481.440 569.665 ;
        RECT 483.840 17.175 558.240 569.665 ;
        RECT 560.640 17.175 573.785 569.665 ;
  END
END coefio
END LIBRARY

